module project_fulltest;

    // Parameters
    localparam wordsize = 32;
    localparam Nreg = 32;
    localparam Nchars = 64;
    localparam charcode_size = $clog2(Nchars);
    localparam bmem_size = Nchars * 256;
    localparam smem_size = 1200;


    // Inputs
    logic clk;
    logic reset;
    logic [wordsize-1:0] keyb_char, accel_val;  // for simulation, directly feed keyb_char and accel_var from tester

     
     
     
    // Signals connected to the instruction memory
    wire [31:0] pc             =uut.pc;                     // PC
    wire [31:0] instr          =uut.instr;                  // instr coming out of instr mem
    
    // Signals connected to the memory + IO unit
    wire [31:0] mem_addr       =uut.mem_addr;               // addr sent to data mem
    wire        wr             =uut.mips.c.wr;              // write enable produced by controller
    wire        mem_wr         =uut.mem_wr;                // write enable reaching inside data mem
    wire [31:0] mem_readdata   =uut.mem_readdata;           // data read from data mem
    wire [31:0] mem_writedata  =uut.mem_writedata;               // write data reaching inside data mem

    // Control inputs/output of the ALU (module uut.mips.dp.alu)
    wire  [4:0] alufn          =uut.mips.dp.alu.ALUfn;      // ALU function
    wire        Z              =uut.mips.Z;                 // Zero flag

    // Data values inside the datapath (module uut.mips.dp)
    wire [31:0] ReadData1      =uut.mips.dp.ReadData1;       // Reg[rs]
    wire [31:0] ReadData2      =uut.mips.dp.ReadData2;       // Reg[rt]
    wire [31:0] alu_result     =uut.mips.dp.alu_result;      // ALU's output
    wire [31:0] signImm        =uut.mips.dp.signImm;         // sign-/zero-extended immediate
    wire [31:0] aluA           =uut.mips.dp.aluA;            // operand A for ALU
    wire [31:0] aluB           =uut.mips.dp.aluB;            // operand B for ALU

    // Updates to the register file (module uut.mips.dp.rf)
    wire        werf           =uut.mips.dp.rf.wr;          // WERF = write enable for register file
    wire [4:0]  reg_writeaddr  =uut.mips.dp.rf.WriteAddr;    // destination register
    wire [31:0] reg_writedata  =uut.mips.dp.rf.WriteData;    // write data for register file

    // Control signals inside the datapath (module uut.mips.dp)
    wire [1:0] pcsel           =uut.mips.dp.pcsel;
    wire [1:0] wasel           =uut.mips.dp.wasel;
    wire sgnext                =uut.mips.dp.sgnext;
    wire bsel                  =uut.mips.dp.bsel;
    wire [1:0] wdsel           =uut.mips.dp.wdsel;
    wire [1:0] asel            =uut.mips.dp.asel;
    
    // Signals related to the memory + IO unit (module memIO)
    wire [$clog2(smem_size)-1:0] smem_addr   =uut.smem_addr;             // address from vgadisplaydriver to access screen mem
    wire [charcode_size-1:0]  charcode       =uut.charcode;              // character code returned by screen mem
    wire cpu_wr                =uut.memIO.cpu_wr;
    wire dmem_wr               =uut.memIO.dmem_wr;
    wire smem_wr               =uut.memIO.smem_wr;
    wire sound_wr              =uut.memIO.sound_wr;
    wire lights_wr             =uut.memIO.lights_wr;
    wire [31:0] smem_readdata  =uut.memIO.smem_readdata;
    wire [31:0] dmem_readdata  =uut.memIO.dmem_readdata;
    wire [31:0] keyb_char      =uut.memIO.keyb_char;
    wire [31:0] accel_val      =uut.memIO.accel_val;
    wire [31:0] cpu_addr       =uut.memIO.cpu_addr;
    wire [31:0] cpu_readdata   =uut.memIO.cpu_readdata;
    wire [31:0] cpu_writedata  =uut.memIO.cpu_writedata;
   
    // Signals related to display driver (module vgadisplaydriver)
    wire hsync                 =uut.hsync;
    wire vsync                 =uut.vsync;
    wire [3:0] red             =uut.red;
    wire [3:0] green           =uut.green;
    wire [3:0] blue            =uut.blue;
    wire [9:0] x               =uut.display.x;
    wire [9:0] y               =uut.display.y;
    wire [$clog2(bmem_size)-1:0] bmem_addr =uut.display.bmem_addr;
    wire [11:0] bmem_color     =uut.display.bmem_color;

    // Other I/O signals (sound and lights) inside top-level module uut
    wire [31:0] period         =uut.period;                // period for sound module
    wire [15:0] LED            =uut.LED;                   // light pattern for LEDs    


    // Instantiate the Unit Under Test (UUT)
    top #(
      .wordsize(wordsize),                // word size for the processor
      .Nreg(Nreg),                        // number of registers
      .Nchars(Nchars),                    // number of characters/sprites
      .imem_size(1024),                   // imem size, must be >= # instructions in program
      .imem_init("imem_fulltest_nopause.mem"),    // program code
      .dmem_size(1024),                   // dmem size, must be >= # words in .data of program + size of stack
      .dmem_init("dmem_test.mem"),        // program data + stack space
      .smem_init("smem_test.mem"), 	      // text file to initialize screen memory
      .bmem_init("bmem_test.mem")         // sprite definitions
    ) uut(
      .clk, .reset,
      .keyb_char, .accel_val  // for simulation, directly feed keyb_char and accel_var from tester
    );

//
// CHECK ALL VALUES ABOVE THIS LINE
// YOU SHOULD NOT NEED TO MODIFY ANYTHING BELOW
//

   initial begin
      // Initialize Inputs
      clk = 0;
      reset = 0;
      keyb_char = 0;
      accel_val = 0;
   end
    
   initial begin    
      #200 keyb_char = 32'h1D;
      #200 keyb_char = 32'h23;
      #200 keyb_char = 32'h1B;
      #200 keyb_char = 32'h1C;
   end
    
   initial begin
      logic [8:0] accelX=0, accelY=0;
      forever begin
         #20
         accelX += 10;
         accelY += 10;
         accel_val = {7'b0, accelX[8:0], 7'b0, accelY[8:0]};
      end
   end

   initial begin
      #0.5 clk = 0;
      forever
         #0.5 clk <= ~clk;
   end
   
   initial begin
      #1000 $finish;
   end
   
   
   
   // SELF-CHECKING CODE
   
   selfcheck_nopause #(.Nchars(Nchars), .smem_size(smem_size)) c();

    wire [31:0] c_pc=c.pc;
    wire [31:0] c_instr=c.instr;
    wire [31:0] c_mem_addr=c.mem_addr;
    wire        c_mem_wr=c.mem_wr;
    wire [31:0] c_mem_readdata=c.mem_readdata;
    wire [31:0] c_mem_writedata=c.mem_writedata;
    wire [31:0] c_period=c.period;
    wire [15:0] c_LED=c.LED;
    wire        c_werf=c.werf;
    wire  [4:0] c_alufn=c.alufn;
    wire        c_Z=c.Z;
    wire [31:0] c_ReadData1=c.ReadData1;
    wire [31:0] c_ReadData2=c.ReadData2;
    wire [31:0] c_alu_result=c.alu_result;
    wire [4:0]  c_reg_writeaddr=c.reg_writeaddr;
    wire [31:0] c_reg_writedata=c.reg_writedata;
    wire [31:0] c_signImm=c.signImm;
    wire [31:0] c_aluA=c.aluA;
    wire [31:0] c_aluB=c.aluB;
    wire [1:0]  c_pcsel=c.pcsel;
    wire [1:0]  c_wasel=c.wasel;
    wire        c_sgnext=c.sgnext;
    wire        c_bsel=c.bsel;
    wire [1:0]  c_wdsel=c.wdsel;
    wire        c_wr=c.wr;
    wire [1:0]  c_asel=c.asel;
    wire [10:0] c_smem_addr=c.smem_addr;
    wire [charcode_size-1:0]  c_charcode=c.charcode;
    wire        c_dmem_wr=c.dmem_wr;
    wire        c_smem_wr=c.smem_wr;
    wire        c_hsync=c.hsync;
    wire        c_vsync=c.vsync;
    wire [3:0]  c_red=c.red;
    wire [3:0]  c_green=c.green;
    wire [3:0]  c_blue=c.blue;
    wire [9:0]  c_x=c.x;
    wire [9:0]  c_y=c.y;
    wire [$clog2(bmem_size)-1:0] c_bmem_addr=c.bmem_addr;
    wire [11:0] c_bmem_color=c.bmem_color;
    wire c_sound_wr=c.sound_wr;
    wire c_lights_wr=c.lights_wr;
    wire [31:0] c_smem_readdata=c.smem_readdata;
    wire [31:0] c_dmem_readdata=c.dmem_readdata;
    wire [31:0] c_keyb_char=c.keyb_char;
    wire [31:0] c_accel_val=c.accel_val;
    wire [31:0] c_cpu_addr=c.cpu_addr;
    wire [31:0] c_cpu_readdata=c.cpu_readdata;
    wire [31:0] c_cpu_writedata=c.cpu_writedata;
  

  
    function mismatch;  // some trickery needed to match two values with don't cares
        input p, q;      // mismatch in a bit position is ignored if q has an 'x' in that bit
        integer p, q;
        mismatch = (((p ^ q) ^ q) !== q);
    endfunction

    wire ERROR;
    wire ERROR_pc             = mismatch(pc, c.pc) ? 1'bx : 1'b0;
    wire ERROR_instr          = mismatch(instr, c.instr) ? 1'bx : 1'b0;
    wire ERROR_mem_addr       = mismatch(mem_addr, c.mem_addr) ? 1'bx : 1'b0;
    wire ERROR_mem_wr         = mismatch(mem_wr, c.mem_wr) ? 1'bx : 1'b0;
    wire ERROR_mem_readdata   = mismatch(mem_readdata, c.mem_readdata) ? 1'bx : 1'b0;
    wire ERROR_mem_writedata  = c.mem_wr & (mismatch(mem_writedata, c.mem_writedata) ? 1'bx : 1'b0);
    wire ERROR_period         = mismatch(period, c.period) ? 1'bx : 1'b0;
    wire ERROR_LED            = mismatch(LED, c.LED) ? 1'bx : 1'b0;
    wire ERROR_werf           = mismatch(werf, c.werf) ? 1'bx : 1'b0;
    wire ERROR_alufn          = mismatch(alufn, c.alufn) ? 1'bx : 1'b0;
    wire ERROR_Z              = mismatch(Z, c.Z) ? 1'bx : 1'b0;
    wire ERROR_ReadData1      = mismatch(ReadData1, c.ReadData1) ? 1'bx : 1'b0;
    wire ERROR_ReadData2      = mismatch(ReadData2, c.ReadData2) ? 1'bx : 1'b0;
    wire ERROR_alu_result     = mismatch(alu_result, c.alu_result) ? 1'bx : 1'b0;
    wire ERROR_reg_writeaddr  = c.werf & (mismatch(reg_writeaddr, c.reg_writeaddr) ? 1'bx : 1'b0);
    wire ERROR_reg_writedata  = c.werf & (mismatch(reg_writedata, c.reg_writedata) ? 1'bx : 1'b0);
    wire ERROR_signImm        = mismatch(signImm, c.signImm) ? 1'bx : 1'b0;
    wire ERROR_aluA           = mismatch(aluA, c.aluA) ? 1'bx : 1'b0;
    wire ERROR_aluB           = mismatch(aluB, c.aluB) ? 1'bx : 1'b0;
    wire ERROR_pcsel          = mismatch(pcsel, c.pcsel) ? 1'bx : 1'b0;
    wire ERROR_wasel          = c.werf & (mismatch(wasel, c.wasel) ? 1'bx : 1'b0);
    wire ERROR_sgnext         = mismatch(sgnext, c.sgnext) ? 1'bx : 1'b0;
    wire ERROR_bsel           = mismatch(bsel, c.bsel) ? 1'bx : 1'b0;
    wire ERROR_wdsel          = mismatch(wdsel, c.wdsel) ? 1'bx : 1'b0;
    wire ERROR_wr             = mismatch(wr, c.wr) ? 1'bx : 1'b0;
    wire ERROR_asel           = mismatch(asel, c.asel) ? 1'bx : 1'b0;
    wire ERROR_smem_addr      = mismatch(smem_addr, c.smem_addr) ? 1'bx : 1'b0;
    wire ERROR_charcode       = mismatch(charcode, c.charcode) ? 1'bx : 1'b0;
    wire ERROR_dmem_wr        = mismatch(dmem_wr, c.dmem_wr) ? 1'bx : 1'b0;
    wire ERROR_smem_wr        = mismatch(smem_wr, c.smem_wr) ? 1'bx : 1'b0;
    wire ERROR_sound_wr       = mismatch(sound_wr, c.sound_wr) ? 1'bx : 1'b0;
    wire ERROR_lights_wr      = mismatch(lights_wr, c.lights_wr) ? 1'bx : 1'b0;
    wire ERROR_smem_readdata  = mismatch(smem_readdata, c.smem_readdata) ? 1'bx : 1'b0;
    wire ERROR_dmem_readdata  = mismatch(dmem_readdata, c.dmem_readdata) ? 1'bx : 1'b0;
    wire ERROR_keyb_char      = mismatch(keyb_char, c.keyb_char) ? 1'bx : 1'b0;
    wire ERROR_accel_val      = mismatch(accel_val, c.accel_val) ? 1'bx : 1'b0;
    wire ERROR_cpu_addr       = mismatch(cpu_addr, c.cpu_addr) ? 1'bx : 1'b0;
    wire ERROR_cpu_readdata   = mismatch(cpu_readdata, c.cpu_readdata) ? 1'bx : 1'b0;
    wire ERROR_cpu_writedata  = mismatch(cpu_writedata, c.cpu_writedata) ? 1'bx : 1'b0;  
    wire ERROR_hsync          = mismatch(hsync, c.hsync) ? 1'bx : 1'b0;
    wire ERROR_vsync          = mismatch(vsync, c.vsync) ? 1'bx : 1'b0;
    wire ERROR_red            = mismatch(red, c.red) ? 1'bx : 1'b0;
    wire ERROR_green          = mismatch(green, c.green) ? 1'bx : 1'b0;
    wire ERROR_blue           = mismatch(blue, c.blue) ? 1'bx : 1'b0;
    wire ERROR_x              = mismatch(x, c.x) ? 1'bx : 1'b0;
    wire ERROR_y              = mismatch(y, c.y) ? 1'bx : 1'b0;
    wire ERROR_bmem_addr      = mismatch(bmem_addr, c.bmem_addr) ? 1'bx : 1'b0;
    wire ERROR_bmem_color     = mismatch(bmem_color, c.bmem_color) ? 1'bx : 1'b0;

    assign ERROR = ERROR_pc | ERROR_instr | ERROR_mem_addr | ERROR_mem_wr | ERROR_mem_readdata 
              | ERROR_mem_writedata | ERROR_period | ERROR_LED | ERROR_werf | ERROR_alufn | ERROR_Z
              | ERROR_ReadData1 | ERROR_ReadData2 | ERROR_alu_result | ERROR_reg_writeaddr
              | ERROR_reg_writedata | ERROR_signImm | ERROR_aluA | ERROR_aluB
              | ERROR_pcsel | ERROR_wasel | ERROR_sgnext | ERROR_bsel | ERROR_wdsel | ERROR_wr | ERROR_asel
              | ERROR_smem_addr | ERROR_charcode | ERROR_dmem_wr | ERROR_smem_wr 
              | ERROR_sound_wr | ERROR_lights_wr | ERROR_smem_readdata | ERROR_dmem_readdata
              | ERROR_keyb_char | ERROR_accel_val | ERROR_cpu_addr | ERROR_cpu_readdata | ERROR_cpu_writedata
              | ERROR_hsync | ERROR_vsync
              | ERROR_red | ERROR_green | ERROR_blue | ERROR_x | ERROR_y | ERROR_bmem_addr | ERROR_bmem_color;


    initial begin
        $monitor("#%02d {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h%h, 32'h%h, 32'h%h, 1'b%b, 32'h%h, 32'h%h, 32'h%h, 16'h%h, 1'b%b, 5'b%b, 1'b%b, 32'h%h, 32'h%h, 32'h%h, 5'h%h, 32'h%h, 32'h%h, 32'h%h, 32'h%h, 2'b%b, 2'b%b, 1'b%b, 1'b%b, 2'b%b, 1'b%b, 2'b%b};",
                  $time, pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel);        
        $monitor("#%02d {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b%b, 1'b%b, 1'b%b, 1'b%b, 4'h%h, 4'h%h, 4'h%h, 10'h%h, 10'h%h, 12'h%h};",
                  $time, dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color);
        $monitor("#%02d {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b%b, 1'b%b, 32'h%h, 32'h%h, 32'h%h, 32'h%h, 32'h%h, 32'h%h, 32'h%h};",
                  $time, sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata);
        $monitor("#%02d smem_addr <= 'h%h;", $time, smem_addr);
        $monitor("#%02d bmem_addr <= 'h%h;", $time, bmem_addr);
        $monitor("#%02d charcode  <= 'h%h;", $time, charcode);
    end
    
endmodule



// CHECKER MODULE

module selfcheck_nopause #(
    parameter Nchars=64,
    parameter smem_size=1200,
    localparam charcode_size=$clog2(Nchars),
    localparam bmem_size=Nchars*256
  )(
  );
    logic  [31:0] pc;
    logic  [31:0] instr;
    logic  [31:0] mem_addr;
    logic         mem_wr;
    logic  [31:0] mem_readdata;
    logic  [31:0] mem_writedata;
    logic  [31:0] period;
    logic  [15:0] LED;
    logic         werf;
    logic   [4:0] alufn;
    logic         Z;
    logic  [31:0] ReadData1;
    logic  [31:0] ReadData2;
    logic  [31:0] alu_result;
    logic  [4:0]  reg_writeaddr;
    logic  [31:0] reg_writedata;
    logic  [31:0] signImm;
    logic  [31:0] aluA;
    logic  [31:0] aluB;
    logic   [1:0] pcsel;
    logic   [1:0] wasel;
    logic         sgnext;
    logic         bsel;
    logic   [1:0] wdsel;
    logic         wr;
    logic   [1:0] asel;
    logic  [$clog2(smem_size)-1:0] smem_addr;
    logic  [charcode_size-1:0] charcode;
    logic dmem_wr;
    logic smem_wr;
    logic hsync;
    logic vsync;
    logic   [3:0] red;
    logic   [3:0] green;
    logic   [3:0] blue;
    logic   [9:0] x;
    logic   [9:0] y;
    logic  [$clog2(bmem_size)-1:0] bmem_addr;
    logic  [11:0] bmem_color;
    logic         sound_wr, lights_wr;
    logic  [31:0] smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata;
    
initial begin
fork

#00 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400000, 32'h3c1d1001, 32'h10010000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h10010000, 5'h1d, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#00 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h000, 10'h000, 12'hf20};
#00 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010000, 32'h00000000, 32'hxxxxxxxx};
#00 smem_addr <= 'h000;
#00 bmem_addr <= 'h0000;
#00 charcode  <= 'h00;
#01 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400004, 32'h37bd1000, 32'h10011000, 1'b0, 32'h00000000, 32'h10010000, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'h10010000, 32'h10011000, 5'h1d, 32'h10011000, 32'h00001000, 32'h10010000, 32'h00001000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#01 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10011000, 32'h00000000, 32'h10010000};
#02 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400008, 32'h23befffc, 32'h10010ffc, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'hxxxxxxxx, 32'h10010ffc, 5'h1e, 32'h10010ffc, 32'hfffffffc, 32'h10011000, 32'hfffffffc, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#02 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h00000000, 32'hxxxxxxxx};
#03 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040000c, 32'h24110014, 32'h00000014, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000014, 5'h11, 32'h00000014, 32'h00000014, 32'h00000000, 32'h00000014, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#03 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h00000000, 32'h00000000, 32'h00000014, 32'hxxxxxxxx, 32'hxxxxxxxx};
#04 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400010, 32'h2412000f, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000000f, 5'h12, 32'h0000000f, 32'h0000000f, 32'h00000000, 32'h0000000f, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#04 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000000, 32'h00000000, 32'h0000000f, 32'hxxxxxxxx, 32'hxxxxxxxx};
#04 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h001, 10'h000, 12'hf20};
#04 bmem_addr <= 'h0001;
#05 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h24040002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#05 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 32'hxxxxxxxx};
#06 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00112821, 32'h00000014, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000014, 32'h00000014, 5'h05, 32'h00000014, 32'h00002821, 32'h00000000, 32'h00000014, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#06 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h00000000, 32'h00000000, 32'h00000014, 32'hxxxxxxxx, 32'h00000014};
#07 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h00123021, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h0000000f, 5'h06, 32'h0000000f, 32'h00003021, 32'h00000000, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#07 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000000, 32'h00000000, 32'h0000000f, 32'hxxxxxxxx, 32'h0000000f};
#08 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h002, 10'h000, 12'hf20};
#08 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h0c10003e, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h00400024, 32'h0000003e, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#08 bmem_addr <= 'h0002;
#08 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'hxxxxxxxx};
#09 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000f8, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'h00000000, 32'h10011000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#09 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000000, 32'h10011000};
#10 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h00000000, 32'h00400024, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#10 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010ffc, 32'h00000000, 32'h00400024};
#10 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h002, 10'h000, 12'hf20};
#11 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010ff8, 32'h00000000, 32'hxxxxxxxx};
#11 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'hafa80008, 32'h10010ff8, 1'b1, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#12 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010ff4, 32'h00000000, 32'hxxxxxxxx};
#12 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'hafa90004, 32'h10010ff4, 1'b1, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#12 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h003, 10'h000, 12'hf20};
#12 bmem_addr <= 'h0003;
#13 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10010ff0, 32'h00000000, 32'hxxxxxxxx};
#13 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#14 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h10020000, 32'h00000000, 32'hxxxxxxxx};
#14 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#14 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h003, 10'h000, 12'hf20};
#15 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'hxxxxxxxx, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#16 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h00064940, 32'h000001e0, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h000001e0, 5'h09, 32'h000001e0, 32'h00004940, 32'h00000005, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#16 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h000001e0, 32'hxxxxxxxx, 32'h0000000f};
#16 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h004, 10'h000, 12'hf20};
#16 bmem_addr <= 'h0004;
#17 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h000650c0, 32'h00000078, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000078, 5'h0a, 32'h00000078, 32'h000050c0, 32'h00000003, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#17 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000078, 32'hxxxxxxxx, 32'h0000000f};
#18 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h012a4820, 32'h00000258, 1'b0, 32'hxxxxxxxx, 32'h00000078, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h000001e0, 32'h00000078, 32'h00000258, 5'h09, 32'h00000258, 32'h00004820, 32'h000001e0, 32'h00000078, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#18 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000258, 32'hxxxxxxxx, 32'h00000078};
#19 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h01254820, 32'h0000026c, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000258, 32'h00000014, 32'h0000026c, 5'h09, 32'h0000026c, 32'h00004820, 32'h00000258, 32'h00000014, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#19 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h0000026c, 32'hxxxxxxxx, 32'h00000014};
#20 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h000a000a, 32'h000009b0, 32'hxxxxxxxx, 32'h0000026c};
#20 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h00094880, 32'h000009b0, 1'b0, 32'hxxxxxxxx, 32'h0000026c, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000026c, 32'h000009b0, 5'h09, 32'h000009b0, 32'h00004880, 32'h00000002, 32'h0000026c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#20 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h005, 10'h000, 12'hf20};
#20 bmem_addr <= 'h0005;
#21 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h01094020, 32'h100209b0, 1'b0, 32'h00000000, 32'h000009b0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000009b0, 32'h100209b0, 5'h08, 32'h100209b0, 32'h00004020, 32'h10020000, 32'h000009b0, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#21 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h000a000a, 32'h100209b0, 32'h00000000, 32'h000009b0};
#22 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'had040000, 32'h100209b0, 1'b1, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h100209b0, 32'h00000002, 32'h100209b0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100209b0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#22 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h000a000a, 32'h100209b0, 32'h00000000, 32'h00000002};
#22 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h005, 10'h000, 12'hf20};
#23 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h00000000, 32'h000a000a, 32'h10010ffc, 32'h00400024, 32'h00400024};
#23 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h00400024, 32'h00400024, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'h1f, 32'h00400024, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#23 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h005, 10'h000, 12'hf20};
#24 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h006, 10'h000, 12'hf20};
#24 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h100209b0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100209b0, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#24 bmem_addr <= 'h0006;
#24 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h000a000a, 32'h10010ff8, 32'hxxxxxxxx, 32'h100209b0};
#25 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h000009b0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000009b0, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#25 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h000a000a, 32'h10010ff4, 32'hxxxxxxxx, 32'h000009b0};
#26 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000078, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000078, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#26 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h000a000a, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000078};
#27 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#27 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h000a000a, 32'h10011000, 32'h00000000, 32'h10010ff0};
#28 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400144, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400024, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#28 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h000a000a, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#28 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h007, 10'h000, 12'hf20};
#28 bmem_addr <= 'h0007;
#29 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h0c1000d3, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h00400028, 32'h000000d3, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#29 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h000a000a, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'hxxxxxxxx};
#30 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040034c, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10020000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#30 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h000a000a, 32'h10030000, 32'h00000000, 32'h10020000};
#31 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400350, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#31 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h000a000a, 32'h10030000, 32'h00000000, 32'h00000000};
#32 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h008, 10'h000, 12'hf20};
#32 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400354, 32'h8c220004, 32'h10030004, 1'b0, 32'h000a000a, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'hxxxxxxxx, 32'h10030004, 5'h02, 32'h000a000a, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#32 bmem_addr <= 'h0008;
#32 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000000, 32'h000a000a, 32'h10030004, 32'h000a000a, 32'hxxxxxxxx};
#33 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400358, 32'h00021402, 32'h0000000a, 1'b0, 32'hxxxxxxxx, 32'h000a000a, 32'h00000000, 16'h0000, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h000a000a, 32'h0000000a, 5'h02, 32'h0000000a, 32'h00001402, 32'h00000010, 32'h000a000a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#33 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000000, 32'h000a000a, 32'h0000000a, 32'hxxxxxxxx, 32'h000a000a};
#34 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040035c, 32'h304201ff, 32'h0000000a, 1'b0, 32'hxxxxxxxx, 32'h0000000a, 32'h00000000, 16'h0000, 1'b1, 5'bx0000, 1'b0, 32'h0000000a, 32'h0000000a, 32'h0000000a, 5'h02, 32'h0000000a, 32'h000001ff, 32'h0000000a, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#34 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000000, 32'h000a000a, 32'h0000000a, 32'hxxxxxxxx, 32'h0000000a};
#35 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400360, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400028, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#35 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h000a000a, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#36 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h009, 10'h000, 12'hf20};
#36 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h00022300, 32'h0000a000, 1'b0, 32'hxxxxxxxx, 32'h0000000a, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000a, 32'h0000a000, 5'h04, 32'h0000a000, 32'h00002300, 32'h0000000c, 32'h0000000a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#36 bmem_addr <= 'h0009;
#36 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h000a000a, 32'h0000a000, 32'hxxxxxxxx, 32'h0000000a};
#37 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h0c1000de, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h00400030, 32'h000000de, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#37 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h000a000a, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'hxxxxxxxx};
#38 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400378, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h00000000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#38 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h000a000a, 32'h10030000, 32'h00000000, 32'h10030000};
#39 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040037c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#39 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h000a000a, 32'h10030000, 32'h00000000, 32'h00000000};
#40 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000000, 32'h00140014, 32'h10030008, 32'hxxxxxxxx, 32'h0000a000};
#40 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h00a, 10'h000, 12'hf20};
#40 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400380, 32'hac240008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h0000a000, 32'h00000000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h0000a000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#40 bmem_addr <= 'h000a;
#41 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400384, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0000a000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400030, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#41 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00140014, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#42 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h0c1000d9, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0000a000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h00400034, 32'h000000d9, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#42 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00140014, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'hxxxxxxxx};
#43 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400364, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h0000a000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#43 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00140014, 32'h10030000, 32'h00000000, 32'h10030000};
#44 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h00b, 10'h000, 12'hf20};
#44 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400368, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h0000a000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#44 bmem_addr <= 'h000b;
#44 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00140014, 32'h10030000, 32'h00000000, 32'h00000000};
#45 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040036c, 32'h8c220004, 32'h10030004, 1'b0, 32'h00140014, 32'h0000000a, 32'h0000a000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h0000000a, 32'h10030004, 5'h02, 32'h00140014, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#45 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000000, 32'h00140014, 32'h10030004, 32'h00140014, 32'h0000000a};
#46 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400370, 32'h304201ff, 32'h00000014, 1'b0, 32'hxxxxxxxx, 32'h00140014, 32'h0000a000, 16'h0000, 1'b1, 5'bx0000, 1'b0, 32'h00140014, 32'h00140014, 32'h00000014, 5'h02, 32'h00000014, 32'h000001ff, 32'h00140014, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#46 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h00000000, 32'h00140014, 32'h00000014, 32'hxxxxxxxx, 32'h00140014};
#47 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400374, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0000a000, 16'h0000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400034, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#47 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00140014, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#48 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h00c, 10'h000, 12'hf20};
#48 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h00021142, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h0000a000, 16'h0000, 1'b1, 5'bx1010, 1'b1, 32'h00000000, 32'h00000014, 32'h00000000, 5'h02, 32'h00000000, 32'h00001142, 32'h00000005, 32'h00000014, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#48 bmem_addr <= 'h000c;
#48 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00140014, 32'h00000000, 32'hxxxxxxxx, 32'h00000014};
#49 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h24040001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h0000a000, 32'h0000a000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000a000, 32'h00000001, 5'h04, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#49 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00140014, 32'h00000001, 32'hxxxxxxxx, 32'h0000a000};
#50 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h00442004, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h0000a000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h00000001, 5'h04, 32'h00000001, 32'h00002004, 32'h00000000, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#50 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00140014, 32'h00000001, 32'hxxxxxxxx, 32'h00000001};
#51 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h0c1000e6, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0000a000, 16'h0000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h00400044, 32'h000000e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#51 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00140014, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'hxxxxxxxx};
#52 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400398, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h0000a000, 16'h0000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#52 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h00d, 10'h000, 12'hf20};
#52 bmem_addr <= 'h000d;
#52 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00140014, 32'h10030000, 32'h00000000, 32'h10030000};
#53 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040039c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h0000a000, 16'h0000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#53 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00140014, 32'h10030000, 32'h00000000, 32'h00000000};
#54 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a0, 32'hac24000c, 32'h1003000c, 1'b1, 32'hxxxxxxxx, 32'h00000001, 32'h0000a000, 16'h0000, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000001, 32'h1003000c, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10030000, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#54 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b1, 32'h00000003, 32'h00000023, 32'h00000000, 32'h00140014, 32'h1003000c, 32'hxxxxxxxx, 32'h00000001};
#55 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a4, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0000a000, 16'h0001, 1'b0, 5'bxxxxx, 1'bx, 32'h00400044, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#55 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00140014, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#56 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h00e, 10'h000, 12'hf20};
#56 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h2404000f, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h0000a000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000001, 32'h0000000f, 5'h04, 32'h0000000f, 32'h0000000f, 32'h00000000, 32'h0000000f, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#56 bmem_addr <= 'h000e;
#56 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000000, 32'h00140014, 32'h0000000f, 32'hxxxxxxxx, 32'h00000001};
#57 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h0c100066, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0000a000, 16'h0001, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'hxxxxxxxx, 32'hxxxxxxxx, 5'h1f, 32'h0040004c, 32'h00000066, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#57 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00140014, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'hxxxxxxxx};
#58 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h0000a000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#58 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00140014, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#59 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h00400024, 32'h0040004c, 32'h0000a000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#59 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h00000000, 32'h00140014, 32'h10010ffc, 32'h00400024, 32'h0040004c};
#59 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h00e, 10'h000, 12'hf20};
#60 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h001e001e, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#60 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0000a000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#60 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h00f, 10'h000, 12'hf20};
#60 bmem_addr <= 'h000f;
#61 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0000a000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#61 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h001e001e, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#62 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0000a000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#62 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h001e001e, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#63 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h0000a000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#63 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h001e001e, 32'h10030000, 32'h00000000, 32'h10030000};
#63 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h00f, 10'h000, 12'hf20};
#64 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h010, 10'h000, 12'h0f0};
#64 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h0000a000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#64 smem_addr <= 'h001;
#64 bmem_addr <= 'h0100;
#64 charcode  <= 'h01;
#64 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h001e001e, 32'h10030000, 32'h00000000, 32'h00000000};
#65 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8c220000, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h0000a000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h02, 32'h00000000, 32'h00000000, 32'h10030000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#66 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h1040000f, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0000a000, 16'h0001, 1'b0, 5'b1xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#66 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h001e001e, 32'h00000000, 32'hxxxxxxxx, 32'h00000000};
#67 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f8, 32'h00021082, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0000a000, 16'h0001, 1'b1, 5'bx1010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h02, 32'h00000000, 32'h00001082, 32'h00000002, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#68 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h011, 10'h000, 12'h0f0};
#68 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001fc, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h0040004c, 32'h0040004c, 32'h0000a000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'h1f, 32'h0040004c, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#68 bmem_addr <= 'h0101;
#68 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h00000000, 32'h001e001e, 32'h10010ffc, 32'h0040004c, 32'h0040004c};
#69 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400200, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0000a000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#69 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h001e001e, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#70 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400204, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0000a000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#70 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h001e001e, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#71 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400208, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0000a000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#71 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h001e001e, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#72 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h012, 10'h000, 12'h0f0};
#72 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040020c, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h0000a000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#72 bmem_addr <= 'h0102;
#72 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h001e001e, 32'h10011000, 32'h00000000, 32'h10010ff0};
#73 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400210, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0000a000, 16'h0001, 1'b0, 5'bxxxxx, 1'bx, 32'h0040004c, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#73 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h001e001e, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#74 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h00028021, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0000a000, 16'h0001, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h10, 32'h00000000, 32'hxxxx8021, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#74 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h001e001e, 32'h00000000, 32'hxxxxxxxx, 32'h00000000};
#75 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h0c1000e2, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0000a000, 16'h0001, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400054, 32'h000000e2, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#75 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h001e001e, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#76 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400388, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h0000a000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#76 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h013, 10'h000, 12'h0f0};
#76 bmem_addr <= 'h0103;
#76 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h001e001e, 32'h10030000, 32'h00000000, 32'h10030000};
#77 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040038c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h0000a000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#77 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h001e001e, 32'h10030000, 32'h00000000, 32'h00000000};
#78 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400390, 32'hac200008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h00000000, 32'h0000a000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#78 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000000, 32'h001e001e, 32'h10030008, 32'hxxxxxxxx, 32'h00000000};
#79 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400394, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0001, 1'b0, 5'bxxxxx, 1'bx, 32'h00400054, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#79 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h001e001e, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#80 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00280028, 32'h00000000, 32'hxxxxxxxx, 32'h00000000};
#80 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h014, 10'h000, 12'h0f0};
#80 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400054, 32'h1200ffef, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0001, 1'b0, 5'b1xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'hffffffef, 32'h00000000, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#80 bmem_addr <= 'h0104;
#81 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h24040002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#81 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00280028, 32'h00000002, 32'hxxxxxxxx, 32'h0000000f};
#82 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00112821, 32'h00000014, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000014, 32'h00000014, 5'h05, 32'h00000014, 32'h00002821, 32'h00000000, 32'h00000014, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#82 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h00000000, 32'h00280028, 32'h00000014, 32'hxxxxxxxx, 32'h00000014};
#83 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h00123021, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h0000000f, 5'h06, 32'h0000000f, 32'h00003021, 32'h00000000, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#83 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000000, 32'h00280028, 32'h0000000f, 32'hxxxxxxxx, 32'h0000000f};
#84 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h015, 10'h000, 12'h0f0};
#84 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h0c10003e, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0001, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400024, 32'h0000003e, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#84 bmem_addr <= 'h0105;
#84 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00280028, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#85 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000f8, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#85 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00280028, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#86 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h0040004c, 32'h00400024, 32'h00000000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#86 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h00000000, 32'h00280028, 32'h10010ffc, 32'h0040004c, 32'h00400024};
#86 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h015, 10'h000, 12'h0f0};
#87 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00280028, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#87 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#88 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h016, 10'h000, 12'h0f0};
#88 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#88 bmem_addr <= 'h0106;
#88 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00280028, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#89 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#89 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00280028, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#90 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'h10030000, 32'h00000000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#90 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00280028, 32'h10020000, 32'h00000000, 32'h10030000};
#90 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h016, 10'h000, 12'h0f0};
#91 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0001, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'hxxxxxxxx, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#91 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00280028, 32'h10020000, 32'h00000000, 32'hxxxxxxxx};
#92 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h00064940, 32'h000001e0, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h000001e0, 5'h09, 32'h000001e0, 32'h00004940, 32'h00000005, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#92 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00280028, 32'h000001e0, 32'hxxxxxxxx, 32'h0000000f};
#92 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h017, 10'h000, 12'h0f0};
#92 bmem_addr <= 'h0107;
#93 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h000650c0, 32'h00000078, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000078, 5'h0a, 32'h00000078, 32'h000050c0, 32'h00000003, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#93 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00280028, 32'h00000078, 32'hxxxxxxxx, 32'h0000000f};
#94 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h012a4820, 32'h00000258, 1'b0, 32'hxxxxxxxx, 32'h00000078, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h000001e0, 32'h00000078, 32'h00000258, 5'h09, 32'h00000258, 32'h00004820, 32'h000001e0, 32'h00000078, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#94 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00280028, 32'h00000258, 32'hxxxxxxxx, 32'h00000078};
#95 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h01254820, 32'h0000026c, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h00000258, 32'h00000014, 32'h0000026c, 5'h09, 32'h0000026c, 32'h00004820, 32'h00000258, 32'h00000014, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#95 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00280028, 32'h0000026c, 32'hxxxxxxxx, 32'h00000014};
#96 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h00094880, 32'h000009b0, 1'b0, 32'hxxxxxxxx, 32'h0000026c, 32'h00000000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000026c, 32'h000009b0, 5'h09, 32'h000009b0, 32'h00004880, 32'h00000002, 32'h0000026c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#96 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 32'h00280028, 32'h000009b0, 32'hxxxxxxxx, 32'h0000026c};
#96 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h018, 10'h000, 12'h0f0};
#96 bmem_addr <= 'h0108;
#97 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h01094020, 32'h100209b0, 1'b0, 32'h00000002, 32'h000009b0, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000009b0, 32'h100209b0, 5'h08, 32'h100209b0, 32'h00004020, 32'h10020000, 32'h000009b0, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#97 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 32'h00280028, 32'h100209b0, 32'h00000002, 32'h000009b0};
#98 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'had040000, 32'h100209b0, 1'b1, 32'h00000002, 32'h00000002, 32'h00000000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h100209b0, 32'h00000002, 32'h100209b0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100209b0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#98 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 32'h00280028, 32'h100209b0, 32'h00000002, 32'h00000002};
#98 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h018, 10'h000, 12'h0f0};
#99 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h00400024, 32'h00400024, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'h1f, 32'h00400024, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#99 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h00000000, 32'h00280028, 32'h10010ffc, 32'h00400024, 32'h00400024};
#99 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h018, 10'h000, 12'h0f0};
#100 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00320032, 32'h10010ff8, 32'hxxxxxxxx, 32'h100209b0};
#100 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h019, 10'h000, 12'h0f0};
#100 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h100209b0, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100209b0, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#100 bmem_addr <= 'h0109;
#101 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h000009b0, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000009b0, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#101 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00320032, 32'h10010ff4, 32'hxxxxxxxx, 32'h000009b0};
#102 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000078, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000078, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#102 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00320032, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000078};
#103 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#103 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00320032, 32'h10011000, 32'h00000000, 32'h10010ff0};
#104 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400144, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0001, 1'b0, 5'bxxxxx, 1'bx, 32'h00400024, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#104 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00320032, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#104 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01a, 10'h000, 12'h0f0};
#104 bmem_addr <= 'h010a;
#105 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h0c1000d3, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0001, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400028, 32'h000000d3, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#106 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040034c, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10020000, 32'h00000000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#106 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00320032, 32'h10030000, 32'h00000000, 32'h10020000};
#107 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400350, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#107 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00320032, 32'h10030000, 32'h00000000, 32'h00000000};
#108 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01b, 10'h000, 12'h0f0};
#108 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400354, 32'h8c220004, 32'h10030004, 1'b0, 32'h00320032, 32'h00000000, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030004, 5'h02, 32'h00320032, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#108 bmem_addr <= 'h010b;
#108 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000000, 32'h00320032, 32'h10030004, 32'h00320032, 32'h00000000};
#109 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400358, 32'h00021402, 32'h00000032, 1'b0, 32'hxxxxxxxx, 32'h00320032, 32'h00000000, 16'h0001, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00320032, 32'h00000032, 5'h02, 32'h00000032, 32'h00001402, 32'h00000010, 32'h00320032, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#109 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 32'h00320032, 32'h00000032, 32'hxxxxxxxx, 32'h00320032};
#110 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040035c, 32'h304201ff, 32'h00000032, 1'b0, 32'hxxxxxxxx, 32'h00000032, 32'h00000000, 16'h0001, 1'b1, 5'bx0000, 1'b0, 32'h00000032, 32'h00000032, 32'h00000032, 5'h02, 32'h00000032, 32'h000001ff, 32'h00000032, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#110 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 32'h00320032, 32'h00000032, 32'hxxxxxxxx, 32'h00000032};
#111 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400360, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0001, 1'b0, 5'bxxxxx, 1'bx, 32'h00400028, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#111 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00320032, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#112 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01c, 10'h000, 12'h0f0};
#112 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h00022300, 32'h00032000, 1'b0, 32'h00000000, 32'h00000032, 32'h00000000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000032, 32'h00032000, 5'h04, 32'h00032000, 32'h00002300, 32'h0000000c, 32'h00000032, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#112 bmem_addr <= 'h010c;
#112 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00320032, 32'h00032000, 32'h00000000, 32'h00000032};
#113 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h0c1000de, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0001, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400030, 32'h000000de, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#113 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00320032, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#114 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400378, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h00000000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#114 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00320032, 32'h10030000, 32'h00000000, 32'h10030000};
#115 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040037c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#115 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00320032, 32'h10030000, 32'h00000000, 32'h00000000};
#116 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01d, 10'h000, 12'h0f0};
#116 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400380, 32'hac240008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h00032000, 32'h00000000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00032000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#116 bmem_addr <= 'h010d;
#116 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000000, 32'h00320032, 32'h10030008, 32'hxxxxxxxx, 32'h00032000};
#117 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400384, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0001, 1'b0, 5'bxxxxx, 1'bx, 32'h00400030, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#117 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00320032, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#118 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h0c1000d9, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0001, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400034, 32'h000000d9, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#119 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400364, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h00032000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#119 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00320032, 32'h10030000, 32'h00000000, 32'h10030000};
#120 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h003c003c, 32'h10030000, 32'h00000000, 32'h00000000};
#120 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01e, 10'h000, 12'h0f0};
#120 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400368, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h00032000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#120 bmem_addr <= 'h010e;
#121 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040036c, 32'h8c220004, 32'h10030004, 1'b0, 32'h003c003c, 32'h00000032, 32'h00032000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000032, 32'h10030004, 5'h02, 32'h003c003c, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#121 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000000, 32'h003c003c, 32'h10030004, 32'h003c003c, 32'h00000032};
#122 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400370, 32'h304201ff, 32'h0000003c, 1'b0, 32'hxxxxxxxx, 32'h003c003c, 32'h00032000, 16'h0001, 1'b1, 5'bx0000, 1'b0, 32'h003c003c, 32'h003c003c, 32'h0000003c, 5'h02, 32'h0000003c, 32'h000001ff, 32'h003c003c, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#122 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h003c003c, 32'h0000003c, 32'hxxxxxxxx, 32'h003c003c};
#123 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400374, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0001, 1'b0, 5'bxxxxx, 1'bx, 32'h00400034, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#123 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h003c003c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#124 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h01f, 10'h000, 12'h0f0};
#124 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h00021142, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h0000003c, 32'h00032000, 16'h0001, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h0000003c, 32'h00000001, 5'h02, 32'h00000001, 32'h00001142, 32'h00000005, 32'h0000003c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#124 bmem_addr <= 'h010f;
#124 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h003c003c, 32'h00000001, 32'hxxxxxxxx, 32'h0000003c};
#125 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h24040001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00032000, 32'h00032000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00032000, 32'h00000001, 5'h04, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#125 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h003c003c, 32'h00000001, 32'hxxxxxxxx, 32'h00032000};
#126 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h00442004, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00032000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000001, 32'h00000001, 32'h00000002, 5'h04, 32'h00000002, 32'h00002004, 32'h00000001, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#126 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h003c003c, 32'h00000002, 32'hxxxxxxxx, 32'h00000001};
#127 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h0c1000e6, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0001, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400044, 32'h000000e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#127 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h003c003c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#128 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400398, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h00032000, 16'h0001, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#128 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h020, 10'h000, 12'hfff};
#128 smem_addr <= 'h002;
#128 bmem_addr <= 'h0200;
#128 charcode  <= 'h02;
#128 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h003c003c, 32'h10030000, 32'h00000000, 32'h10030000};
#129 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040039c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h00032000, 16'h0001, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#129 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h003c003c, 32'h10030000, 32'h00000000, 32'h00000000};
#130 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a0, 32'hac24000c, 32'h1003000c, 1'b1, 32'hxxxxxxxx, 32'h00000002, 32'h00032000, 16'h0001, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000002, 32'h1003000c, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10030000, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#130 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b1, 32'h00000003, 32'h00000023, 32'h00000000, 32'h003c003c, 32'h1003000c, 32'hxxxxxxxx, 32'h00000002};
#131 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a4, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0002, 1'b0, 5'bxxxxx, 1'bx, 32'h00400044, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#131 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h003c003c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#132 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h021, 10'h000, 12'hfff};
#132 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h2404000f, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00032000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h0000000f, 5'h04, 32'h0000000f, 32'h0000000f, 32'h00000000, 32'h0000000f, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#132 bmem_addr <= 'h0201;
#132 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000000, 32'h003c003c, 32'h0000000f, 32'hxxxxxxxx, 32'h00000002};
#133 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h0c100066, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0002, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h0040004c, 32'h00000066, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#133 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h003c003c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#134 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00032000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#134 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h003c003c, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#135 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h00400024, 32'h0040004c, 32'h00032000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#135 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h00000000, 32'h003c003c, 32'h10010ffc, 32'h00400024, 32'h0040004c};
#135 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h021, 10'h000, 12'hfff};
#136 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h003c003c, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#136 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00032000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#136 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h022, 10'h000, 12'hfff};
#136 bmem_addr <= 'h0202;
#137 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00032000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#137 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h003c003c, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#138 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00032000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#138 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h003c003c, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#139 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h00032000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#139 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h003c003c, 32'h10030000, 32'h00000000, 32'h10030000};
#139 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h022, 10'h000, 12'hfff};
#140 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00460046, 32'h10030000, 32'h00000000, 32'h00000000};
#140 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h023, 10'h000, 12'hfff};
#140 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h00032000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#140 bmem_addr <= 'h0203;
#141 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8c220000, 32'h10030000, 1'b0, 32'h00000000, 32'h00000001, 32'h00032000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000001, 32'h10030000, 5'h02, 32'h00000000, 32'h00000000, 32'h10030000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#141 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00460046, 32'h10030000, 32'h00000000, 32'h00000001};
#142 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h1040000f, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0002, 1'b0, 5'b1xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#142 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00460046, 32'h00000000, 32'hxxxxxxxx, 32'h00000000};
#143 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f8, 32'h00021082, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0002, 1'b1, 5'bx1010, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h02, 32'h00000000, 32'h00001082, 32'h00000002, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#144 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hd, 4'hc, 10'h024, 10'h000, 12'hfdc};
#144 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001fc, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h0040004c, 32'h0040004c, 32'h00032000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'h1f, 32'h0040004c, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#144 bmem_addr <= 'h0204;
#144 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h00000000, 32'h00460046, 32'h10010ffc, 32'h0040004c, 32'h0040004c};
#145 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400200, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00032000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#145 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00460046, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#146 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400204, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00032000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#146 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00460046, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#147 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400208, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00032000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#147 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00460046, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#148 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h8, 10'h025, 10'h000, 12'hfc8};
#148 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040020c, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00032000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#148 bmem_addr <= 'h0205;
#148 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00460046, 32'h10011000, 32'h00000000, 32'h10010ff0};
#149 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400210, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0002, 1'b0, 5'bxxxxx, 1'bx, 32'h0040004c, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#149 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00460046, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#150 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h00028021, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0002, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'h10, 32'h00000000, 32'hxxxx8021, 32'h00000000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#150 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00460046, 32'h00000000, 32'hxxxxxxxx, 32'h00000000};
#151 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h0c1000e2, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0002, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400054, 32'h000000e2, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#151 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00460046, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#152 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400388, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h00032000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#152 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h026, 10'h000, 12'hfc6};
#152 bmem_addr <= 'h0206;
#152 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00460046, 32'h10030000, 32'h00000000, 32'h10030000};
#153 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040038c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h00032000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#153 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00460046, 32'h10030000, 32'h00000000, 32'h00000000};
#154 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400390, 32'hac200008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h00000000, 32'h00032000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#154 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000000, 32'h00460046, 32'h10030008, 32'hxxxxxxxx, 32'h00000000};
#155 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400394, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0002, 1'b0, 5'bxxxxx, 1'bx, 32'h00400054, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#155 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00460046, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#156 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h027, 10'h000, 12'hfc6};
#156 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400054, 32'h1200ffef, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0002, 1'b0, 5'b1xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'hffffffef, 32'h00000000, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#156 bmem_addr <= 'h0207;
#156 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00460046, 32'h00000000, 32'hxxxxxxxx, 32'h00000000};
#157 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h24040002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#157 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00460046, 32'h00000002, 32'hxxxxxxxx, 32'h0000000f};
#158 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00112821, 32'h00000014, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000014, 32'h00000014, 5'h05, 32'h00000014, 32'h00002821, 32'h00000000, 32'h00000014, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#158 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h00000000, 32'h00460046, 32'h00000014, 32'hxxxxxxxx, 32'h00000014};
#159 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h00123021, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h0000000f, 5'h06, 32'h0000000f, 32'h00003021, 32'h00000000, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#159 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000000, 32'h00460046, 32'h0000000f, 32'hxxxxxxxx, 32'h0000000f};
#160 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h00500050, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#160 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h028, 10'h000, 12'hfc6};
#160 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h0c10003e, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0002, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400024, 32'h0000003e, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#160 bmem_addr <= 'h0208;
#161 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000f8, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#161 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00500050, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#162 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h0040004c, 32'h00400024, 32'h00000000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#162 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h00000000, 32'h00500050, 32'h10010ffc, 32'h0040004c, 32'h00400024};
#162 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h028, 10'h000, 12'hfc6};
#163 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00500050, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#163 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#164 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h029, 10'h000, 12'hfc6};
#164 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#164 bmem_addr <= 'h0209;
#164 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00500050, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#165 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#165 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00500050, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#166 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'h10030000, 32'h00000000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#166 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00500050, 32'h10020000, 32'h00000000, 32'h10030000};
#166 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h029, 10'h000, 12'hfc6};
#167 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0002, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'hxxxxxxxx, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#167 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00500050, 32'h10020000, 32'h00000000, 32'hxxxxxxxx};
#168 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h00064940, 32'h000001e0, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h000001e0, 5'h09, 32'h000001e0, 32'h00004940, 32'h00000005, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#168 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00500050, 32'h000001e0, 32'hxxxxxxxx, 32'h0000000f};
#168 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h8, 10'h02a, 10'h000, 12'hfc8};
#168 bmem_addr <= 'h020a;
#169 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h000650c0, 32'h00000078, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000078, 5'h0a, 32'h00000078, 32'h000050c0, 32'h00000003, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#169 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00500050, 32'h00000078, 32'hxxxxxxxx, 32'h0000000f};
#170 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h012a4820, 32'h00000258, 1'b0, 32'hxxxxxxxx, 32'h00000078, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h000001e0, 32'h00000078, 32'h00000258, 5'h09, 32'h00000258, 32'h00004820, 32'h000001e0, 32'h00000078, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#170 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00500050, 32'h00000258, 32'hxxxxxxxx, 32'h00000078};
#171 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h01254820, 32'h0000026c, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h00000258, 32'h00000014, 32'h0000026c, 5'h09, 32'h0000026c, 32'h00004820, 32'h00000258, 32'h00000014, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#171 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00500050, 32'h0000026c, 32'hxxxxxxxx, 32'h00000014};
#172 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h00094880, 32'h000009b0, 1'b0, 32'hxxxxxxxx, 32'h0000026c, 32'h00000000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000026c, 32'h000009b0, 5'h09, 32'h000009b0, 32'h00004880, 32'h00000002, 32'h0000026c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#172 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 32'h00500050, 32'h000009b0, 32'hxxxxxxxx, 32'h0000026c};
#172 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'he, 4'hc, 10'h02b, 10'h000, 12'hfec};
#172 bmem_addr <= 'h020b;
#173 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h01094020, 32'h100209b0, 1'b0, 32'h00000002, 32'h000009b0, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000009b0, 32'h100209b0, 5'h08, 32'h100209b0, 32'h00004020, 32'h10020000, 32'h000009b0, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#173 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 32'h00500050, 32'h100209b0, 32'h00000002, 32'h000009b0};
#174 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'had040000, 32'h100209b0, 1'b1, 32'h00000002, 32'h00000002, 32'h00000000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h100209b0, 32'h00000002, 32'h100209b0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100209b0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#174 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 32'h00500050, 32'h100209b0, 32'h00000002, 32'h00000002};
#174 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'he, 4'hc, 10'h02b, 10'h000, 12'hfec};
#175 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h00400024, 32'h00400024, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'h1f, 32'h00400024, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#175 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h00000000, 32'h00500050, 32'h10010ffc, 32'h00400024, 32'h00400024};
#175 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'he, 4'hc, 10'h02b, 10'h000, 12'hfec};
#176 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h02c, 10'h000, 12'hfff};
#176 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h100209b0, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100209b0, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#176 bmem_addr <= 'h020c;
#176 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00500050, 32'h10010ff8, 32'hxxxxxxxx, 32'h100209b0};
#177 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h000009b0, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000009b0, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#177 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00500050, 32'h10010ff4, 32'hxxxxxxxx, 32'h000009b0};
#178 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000078, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000078, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#178 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 32'h00500050, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000078};
#179 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#179 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00500050, 32'h10011000, 32'h00000000, 32'h10010ff0};
#180 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h005a005a, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#180 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400144, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0002, 1'b0, 5'bxxxxx, 1'bx, 32'h00400024, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#180 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h02d, 10'h000, 12'hfff};
#180 bmem_addr <= 'h020d;
#181 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h0c1000d3, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0002, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400028, 32'h000000d3, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#182 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040034c, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10020000, 32'h00000000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#182 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h005a005a, 32'h10030000, 32'h00000000, 32'h10020000};
#183 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400350, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#183 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h005a005a, 32'h10030000, 32'h00000000, 32'h00000000};
#184 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h02e, 10'h000, 12'hfff};
#184 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400354, 32'h8c220004, 32'h10030004, 1'b0, 32'h005a005a, 32'h00000000, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030004, 5'h02, 32'h005a005a, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#184 bmem_addr <= 'h020e;
#184 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000000, 32'h005a005a, 32'h10030004, 32'h005a005a, 32'h00000000};
#185 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400358, 32'h00021402, 32'h0000005a, 1'b0, 32'hxxxxxxxx, 32'h005a005a, 32'h00000000, 16'h0002, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h005a005a, 32'h0000005a, 5'h02, 32'h0000005a, 32'h00001402, 32'h00000010, 32'h005a005a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#185 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 32'h005a005a, 32'h0000005a, 32'hxxxxxxxx, 32'h005a005a};
#186 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040035c, 32'h304201ff, 32'h0000005a, 1'b0, 32'hxxxxxxxx, 32'h0000005a, 32'h00000000, 16'h0002, 1'b1, 5'bx0000, 1'b0, 32'h0000005a, 32'h0000005a, 32'h0000005a, 5'h02, 32'h0000005a, 32'h000001ff, 32'h0000005a, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#186 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 32'h005a005a, 32'h0000005a, 32'hxxxxxxxx, 32'h0000005a};
#187 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400360, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0002, 1'b0, 5'bxxxxx, 1'bx, 32'h00400028, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#187 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h005a005a, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#188 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h02f, 10'h000, 12'hfff};
#188 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h00022300, 32'h0005a000, 1'b0, 32'h00000000, 32'h0000005a, 32'h00000000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000005a, 32'h0005a000, 5'h04, 32'h0005a000, 32'h00002300, 32'h0000000c, 32'h0000005a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#188 bmem_addr <= 'h020f;
#188 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h005a005a, 32'h0005a000, 32'h00000000, 32'h0000005a};
#189 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h0c1000de, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0002, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400030, 32'h000000de, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#189 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h005a005a, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#190 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400378, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h00000000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#190 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h005a005a, 32'h10030000, 32'h00000000, 32'h10030000};
#191 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040037c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#191 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h005a005a, 32'h10030000, 32'h00000000, 32'h00000000};
#192 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h030, 10'h000, 12'hccc};
#192 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400380, 32'hac240008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h0005a000, 32'h00000000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h0005a000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#192 smem_addr <= 'h003;
#192 bmem_addr <= 'h0300;
#192 charcode  <= 'h03;
#192 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000000, 32'h005a005a, 32'h10030008, 32'hxxxxxxxx, 32'h0005a000};
#193 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400384, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0002, 1'b0, 5'bxxxxx, 1'bx, 32'h00400030, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#193 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h005a005a, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#194 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h0c1000d9, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0002, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400034, 32'h000000d9, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#195 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400364, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000000, 32'h10030000, 32'h0005a000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#195 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h005a005a, 32'h10030000, 32'h00000000, 32'h10030000};
#196 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h031, 10'h000, 12'hccc};
#196 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400368, 32'h00200821, 32'h10030000, 1'b0, 32'h00000000, 32'h00000000, 32'h0005a000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#196 bmem_addr <= 'h0301;
#196 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 32'h005a005a, 32'h10030000, 32'h00000000, 32'h00000000};
#197 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040036c, 32'h8c220004, 32'h10030004, 1'b0, 32'h005a005a, 32'h0000005a, 32'h0005a000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h0000005a, 32'h10030004, 5'h02, 32'h005a005a, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#197 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000000, 32'h005a005a, 32'h10030004, 32'h005a005a, 32'h0000005a};
#198 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400370, 32'h304201ff, 32'h0000005a, 1'b0, 32'hxxxxxxxx, 32'h005a005a, 32'h0005a000, 16'h0002, 1'b1, 5'bx0000, 1'b0, 32'h005a005a, 32'h005a005a, 32'h0000005a, 5'h02, 32'h0000005a, 32'h000001ff, 32'h005a005a, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#198 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000000, 32'h005a005a, 32'h0000005a, 32'hxxxxxxxx, 32'h005a005a};
#199 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400374, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0002, 1'b0, 5'bxxxxx, 1'bx, 32'h00400034, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#199 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000000, 32'h005a005a, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#200 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00640064, 32'h00000002, 32'hxxxxxxxx, 32'h0000005a};
#200 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h032, 10'h000, 12'hccc};
#200 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h00021142, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000005a, 32'h0005a000, 16'h0002, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h0000005a, 32'h00000002, 5'h02, 32'h00000002, 32'h00001142, 32'h00000005, 32'h0000005a, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#200 bmem_addr <= 'h0302;
#201 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h24040001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h0005a000, 32'h0005a000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0005a000, 32'h00000001, 5'h04, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#201 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00640064, 32'h00000001, 32'hxxxxxxxx, 32'h0005a000};
#202 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h00442004, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h0005a000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000002, 32'h00000001, 32'h00000004, 5'h04, 32'h00000004, 32'h00002004, 32'h00000002, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#202 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001d, 32'h00640064, 32'h00000004, 32'hxxxxxxxx, 32'h00000001};
#203 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h0c1000e6, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0002, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h00400044, 32'h000000e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#203 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00640064, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#204 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400398, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001d, 32'h10030000, 32'h0005a000, 16'h0002, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#204 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h033, 10'h000, 12'hccc};
#204 bmem_addr <= 'h0303;
#204 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00640064, 32'h10030000, 32'h0000001d, 32'h10030000};
#205 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040039c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001d, 32'h00000000, 32'h0005a000, 16'h0002, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#205 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00640064, 32'h10030000, 32'h0000001d, 32'h00000000};
#206 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a0, 32'hac24000c, 32'h1003000c, 1'b1, 32'hxxxxxxxx, 32'h00000004, 32'h0005a000, 16'h0002, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000004, 32'h1003000c, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10030000, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#206 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b1, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h00640064, 32'h1003000c, 32'hxxxxxxxx, 32'h00000004};
#207 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a4, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0004, 1'b0, 5'bxxxxx, 1'bx, 32'h00400044, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#207 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00640064, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#208 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h034, 10'h000, 12'h999};
#208 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h2404000f, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000004, 32'h0000000f, 5'h04, 32'h0000000f, 32'h0000000f, 32'h00000000, 32'h0000000f, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#208 bmem_addr <= 'h0304;
#208 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h00640064, 32'h0000000f, 32'hxxxxxxxx, 32'h00000004};
#209 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h0c100066, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0004, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000000, 32'hxxxxxxxx, 5'h1f, 32'h0040004c, 32'h00000066, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#209 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00640064, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#210 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#210 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00640064, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#211 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h00400024, 32'h0040004c, 32'h0005a000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#211 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001d, 32'h00640064, 32'h10010ffc, 32'h00400024, 32'h0040004c};
#211 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h034, 10'h000, 12'h999};
#212 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00640064, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#212 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0005a000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#212 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h035, 10'h000, 12'h999};
#212 bmem_addr <= 'h0305;
#213 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0005a000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#213 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00640064, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#214 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0005a000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#214 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00640064, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#215 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001d, 32'h10030000, 32'h0005a000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#215 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00640064, 32'h10030000, 32'h0000001d, 32'h10030000};
#215 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h035, 10'h000, 12'h999};
#216 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h036, 10'h000, 12'h999};
#216 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001d, 32'h00000000, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#216 bmem_addr <= 'h0306;
#216 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00640064, 32'h10030000, 32'h0000001d, 32'h00000000};
#217 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8c220000, 32'h10030000, 1'b0, 32'h0000001d, 32'h00000002, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000002, 32'h10030000, 5'h02, 32'h0000001d, 32'h00000000, 32'h10030000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#217 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00640064, 32'h10030000, 32'h0000001d, 32'h00000002};
#218 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h1040000f, 32'h0000001d, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0004, 1'b0, 5'b1xx01, 1'b0, 32'h0000001d, 32'h00000000, 32'h0000001d, 5'hxx, 32'hxxxxxxxx, 32'h0000000f, 32'h0000001d, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#218 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000004b, 32'h0000001d, 32'h00640064, 32'h0000001d, 32'hxxxxxxxx, 32'h00000000};
#219 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h00024821, 32'h0000001d, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001d, 5'h09, 32'h0000001d, 32'h00004821, 32'h00000000, 32'h0000001d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#219 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000004b, 32'h0000001d, 32'h00640064, 32'h0000001d, 32'hxxxxxxxx, 32'h0000001d};
#220 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h006e006e, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d};
#220 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h037, 10'h000, 12'hf20};
#220 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c0, 32'h24020000, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h0000001d, 32'h00000000, 5'h02, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#220 bmem_addr <= 'h0307;
#221 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c4, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10030000, 32'h0005a000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#221 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h006e006e, 32'h10010000, 32'h00000000, 32'h10030000};
#222 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c8, 32'h34280008, 32'h10010008, 1'b0, 32'h0000001c, 32'hxxxxxxxx, 32'h0005a000, 16'h0004, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010008, 5'h08, 32'h10010008, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#222 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001d, 32'h006e006e, 32'h10010008, 32'h0000001c, 32'hxxxxxxxx};
#223 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001cc, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h0005a000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#223 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h006e006e, 32'h10010000, 32'h00000000, 32'h10010000};
#224 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h038, 10'h000, 12'hf20};
#224 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d0, 32'h342a0018, 32'h10010018, 1'b0, 32'h0000003b, 32'hxxxxxxxx, 32'h0005a000, 16'h0004, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010018, 5'h0a, 32'h10010018, 32'h00000018, 32'h10010000, 32'h00000018, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#224 bmem_addr <= 'h0308;
#224 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h0000001d, 32'h006e006e, 32'h10010018, 32'h0000003b, 32'hxxxxxxxx};
#225 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d4, 32'h01485022, 32'h00000010, 1'b0, 32'hxxxxxxxx, 32'h10010008, 32'h0005a000, 16'h0004, 1'b1, 5'b1xx01, 1'b0, 32'h10010018, 32'h10010008, 32'h00000010, 5'h0a, 32'h00000010, 32'h00005022, 32'h10010018, 32'h10010008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#225 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001d, 32'h006e006e, 32'h00000010, 32'hxxxxxxxx, 32'h10010008};
#226 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h0005a000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#226 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h006e006e, 32'h10010000, 32'h00000000, 32'h10010000};
#227 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#227 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h006e006e, 32'h10010000, 32'h00000000, 32'h00000000};
#228 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h039, 10'h000, 12'hf20};
#228 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010008, 1'b0, 32'h0000001c, 32'h10010008, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h10010008, 32'h10010008, 5'h08, 32'h0000001c, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#228 bmem_addr <= 'h0309;
#228 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001d, 32'h006e006e, 32'h10010008, 32'h0000001c, 32'h10010008};
#229 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000004, 5'h02, 32'h00000004, 32'h00000004, 32'h00000000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#229 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001d, 32'h006e006e, 32'h00000004, 32'hxxxxxxxx, 32'h00000000};
#230 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'hffffffff, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0005a000, 16'h0004, 1'b0, 5'b1xx01, 1'b0, 32'h0000001c, 32'h0000001d, 32'hffffffff, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001c, 32'h0000001d, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#230 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001d, 32'h006e006e, 32'hffffffff, 32'hxxxxxxxx, 32'h0000001d};
#231 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0005a000, 16'h0004, 1'b1, 5'b1x011, 1'b0, 32'h00000004, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h00000004, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#231 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h006e006e, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#232 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h03a, 10'h000, 12'hf20};
#232 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0004, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#232 bmem_addr <= 'h030a;
#232 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h006e006e, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#233 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h0005a000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#233 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h006e006e, 32'h10010000, 32'h00000000, 32'h00000001};
#234 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010004, 1'b0, 32'h00000003, 32'h00000004, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000004, 32'h10010004, 5'h01, 32'h10010004, 32'h00000821, 32'h10010000, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#234 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001d, 32'h006e006e, 32'h10010004, 32'h00000003, 32'h00000004};
#235 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h1001000c, 1'b0, 32'h00000023, 32'h0000001c, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010004, 32'h0000001c, 32'h1001000c, 5'h08, 32'h00000023, 32'h00000008, 32'h10010004, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#235 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h006e006e, 32'h1001000c, 32'h00000023, 32'h0000001c};
#236 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000008, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000004, 32'h00000004, 32'h00000008, 5'h02, 32'h00000008, 32'h00000004, 32'h00000004, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#236 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001d, 32'h006e006e, 32'h00000008, 32'hxxxxxxxx, 32'h00000004};
#236 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h03b, 10'h000, 12'hf20};
#236 bmem_addr <= 'h030b;
#237 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000006, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0005a000, 16'h0004, 1'b0, 5'b1xx01, 1'b0, 32'h00000023, 32'h0000001d, 32'h00000006, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h00000023, 32'h0000001d, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#237 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001d, 32'h006e006e, 32'h00000006, 32'hxxxxxxxx, 32'h0000001d};
#238 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0005a000, 16'h0004, 1'b1, 5'b1x011, 1'b0, 32'h00000008, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h00000008, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#238 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h006e006e, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#239 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0004, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#239 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h006e006e, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#240 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00780078, 32'h10010000, 32'h00000000, 32'h00000001};
#240 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h03c, 10'h000, 12'hf20};
#240 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h0005a000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#240 bmem_addr <= 'h030c;
#241 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010008, 1'b0, 32'h0000001c, 32'h00000008, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000008, 32'h10010008, 5'h01, 32'h10010008, 32'h00000821, 32'h10010000, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#241 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001d, 32'h00780078, 32'h10010008, 32'h0000001c, 32'h00000008};
#242 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010010, 1'b0, 32'h0000001d, 32'h00000023, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010008, 32'h00000023, 32'h10010010, 5'h08, 32'h0000001d, 32'h00000008, 32'h10010008, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#242 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001d, 32'h00780078, 32'h10010010, 32'h0000001d, 32'h00000023};
#243 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h0000000c, 1'b0, 32'hxxxxxxxx, 32'h00000008, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000008, 32'h00000008, 32'h0000000c, 5'h02, 32'h0000000c, 32'h00000004, 32'h00000008, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#243 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h00780078, 32'h0000000c, 32'hxxxxxxxx, 32'h00000008};
#244 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0005a000, 16'h0004, 1'b0, 5'b1xx01, 1'b1, 32'h0000001d, 32'h0000001d, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001d, 32'h0000001d, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#244 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00780078, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d};
#244 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h03d, 10'h000, 12'hf20};
#244 bmem_addr <= 'h030d;
#245 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f8, 32'h00021082, 32'h00000003, 1'b0, 32'hxxxxxxxx, 32'h0000000c, 32'h0005a000, 16'h0004, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000003, 5'h02, 32'h00000003, 32'h00001082, 32'h00000002, 32'h0000000c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#245 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00780078, 32'h00000003, 32'hxxxxxxxx, 32'h0000000c};
#246 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001fc, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h0040004c, 32'h0040004c, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'h1f, 32'h0040004c, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#246 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h0000001d, 32'h00780078, 32'h10010ffc, 32'h0040004c, 32'h0040004c};
#247 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400200, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001d, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#247 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00780078, 32'h10010ff8, 32'hxxxxxxxx, 32'h0000001d};
#248 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400204, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001d, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#248 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00780078, 32'h10010ff4, 32'hxxxxxxxx, 32'h0000001d};
#248 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h03e, 10'h000, 12'hf20};
#248 bmem_addr <= 'h030e;
#249 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400208, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000010, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#249 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00780078, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000010};
#250 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040020c, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#250 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00780078, 32'h10011000, 32'h00000000, 32'h10010ff0};
#251 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400210, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0004, 1'b0, 5'bxxxxx, 1'bx, 32'h0040004c, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#251 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00780078, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#252 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h03f, 10'h000, 12'hf20};
#252 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h00028021, 32'h00000003, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000003, 5'h10, 32'h00000003, 32'hxxxx8021, 32'h00000000, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#252 bmem_addr <= 'h030f;
#252 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00780078, 32'h00000003, 32'hxxxxxxxx, 32'h00000003};
#253 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h0c1000e2, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h0005a000, 16'h0004, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400054, 32'h000000e2, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#253 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00780078, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#254 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400388, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001d, 32'h10010008, 32'h0005a000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010008, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#254 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00780078, 32'h10030000, 32'h0000001d, 32'h10010008};
#255 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040038c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001d, 32'h00000000, 32'h0005a000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#255 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00780078, 32'h10030000, 32'h0000001d, 32'h00000000};
#256 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h040, 10'h000, 12'hf20};
#256 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400390, 32'hac200008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h00000000, 32'h0005a000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#256 smem_addr <= 'h004;
#256 bmem_addr <= 'h0000;
#256 charcode  <= 'h00;
#256 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001d, 32'h00780078, 32'h10030008, 32'hxxxxxxxx, 32'h00000000};
#257 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400394, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0004, 1'b0, 5'bxxxxx, 1'bx, 32'h00400054, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#257 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00780078, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#258 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400054, 32'h1200ffef, 32'h00000003, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0004, 1'b0, 5'b1xx01, 1'b0, 32'h00000003, 32'h00000000, 32'h00000003, 5'hxx, 32'hxxxxxxxx, 32'hffffffef, 32'h00000003, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#258 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00780078, 32'h00000003, 32'hxxxxxxxx, 32'h00000000};
#259 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400058, 32'h20010001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h10030000, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h10030000, 32'h00000001, 5'h01, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#259 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00780078, 32'h00000001, 32'hxxxxxxxx, 32'h10030000};
#260 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001d, 32'h00820082, 32'hfffffffe, 32'hxxxxxxxx, 32'h00000003};
#260 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040005c, 32'h14300005, 32'hfffffffe, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0004, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000003, 32'hfffffffe, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000001, 32'h00000003, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#260 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h041, 10'h000, 12'hf20};
#260 bmem_addr <= 'h0001;
#261 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400074, 32'h20010002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000001, 32'h00000002, 5'h01, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#261 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00820082, 32'h00000002, 32'hxxxxxxxx, 32'h00000001};
#262 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400078, 32'h14300005, 32'hffffffff, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0004, 1'b0, 5'b1xx01, 1'b0, 32'h00000002, 32'h00000003, 32'hffffffff, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000002, 32'h00000003, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#262 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001d, 32'h00820082, 32'hffffffff, 32'hxxxxxxxx, 32'h00000003};
#263 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400090, 32'h20010003, 32'h00000003, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000003, 5'h01, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#263 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00820082, 32'h00000003, 32'hxxxxxxxx, 32'h00000002};
#264 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400094, 32'h14300005, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0004, 1'b0, 5'b1xx01, 1'b1, 32'h00000003, 32'h00000003, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000003, 32'h00000003, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#264 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00820082, 32'h00000000, 32'hxxxxxxxx, 32'h00000003};
#264 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h042, 10'h000, 12'hf20};
#264 bmem_addr <= 'h0002;
#265 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400098, 32'h2252ffff, 32'h0000000e, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h0000000f, 32'h0000000f, 32'h0000000e, 5'h12, 32'h0000000e, 32'hffffffff, 32'h0000000f, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#265 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h00820082, 32'h0000000e, 32'hxxxxxxxx, 32'h0000000f};
#266 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040009c, 32'h0240082a, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0004, 1'b1, 5'b1x011, 1'b1, 32'h0000000e, 32'h00000000, 32'h00000000, 5'h01, 32'h00000000, 32'h0000082a, 32'h0000000e, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#266 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00820082, 32'h00000000, 32'hxxxxxxxx, 32'h00000000};
#267 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000a0, 32'h1020ffdc, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0004, 1'b0, 5'b1xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'hffffffdc, 32'h00000000, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#268 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h043, 10'h000, 12'hf20};
#268 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h24040002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#268 bmem_addr <= 'h0003;
#268 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00820082, 32'h00000002, 32'hxxxxxxxx, 32'h0000000f};
#269 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00112821, 32'h00000014, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000014, 32'h00000014, 5'h05, 32'h00000014, 32'h00002821, 32'h00000000, 32'h00000014, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#269 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h0000001d, 32'h00820082, 32'h00000014, 32'hxxxxxxxx, 32'h00000014};
#270 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h00123021, 32'h0000000e, 1'b0, 32'hxxxxxxxx, 32'h0000000e, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000e, 32'h0000000e, 5'h06, 32'h0000000e, 32'h00003021, 32'h00000000, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#270 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h00820082, 32'h0000000e, 32'hxxxxxxxx, 32'h0000000e};
#271 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h0c10003e, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0004, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400024, 32'h0000003e, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#271 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00820082, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#272 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000f8, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#272 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h044, 10'h000, 12'hf20};
#272 bmem_addr <= 'h0004;
#272 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00820082, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#273 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h0040004c, 32'h00400024, 32'h00000000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#273 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h0000001d, 32'h00820082, 32'h10010ffc, 32'h0040004c, 32'h00400024};
#273 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h044, 10'h000, 12'hf20};
#274 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00820082, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#274 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#275 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#275 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00820082, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#276 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h045, 10'h000, 12'hf20};
#276 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#276 bmem_addr <= 'h0005;
#276 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00820082, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#277 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#277 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00820082, 32'h10020000, 32'h00000000, 32'h00000000};
#277 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h045, 10'h000, 12'hf20};
#278 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0004, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'hxxxxxxxx, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#278 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00820082, 32'h10020000, 32'h00000000, 32'hxxxxxxxx};
#279 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h00064940, 32'h000001c0, 1'b0, 32'hxxxxxxxx, 32'h0000000e, 32'h00000000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000e, 32'h000001c0, 5'h09, 32'h000001c0, 32'h00004940, 32'h00000005, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#279 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00820082, 32'h000001c0, 32'hxxxxxxxx, 32'h0000000e};
#280 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h00000070, 32'hxxxxxxxx, 32'h0000000e};
#280 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h046, 10'h000, 12'hf20};
#280 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h000650c0, 32'h00000070, 1'b0, 32'hxxxxxxxx, 32'h0000000e, 32'h00000000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000070, 5'h0a, 32'h00000070, 32'h000050c0, 32'h00000003, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#280 bmem_addr <= 'h0006;
#281 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h012a4820, 32'h00000230, 1'b0, 32'hxxxxxxxx, 32'h00000070, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h000001c0, 32'h00000070, 32'h00000230, 5'h09, 32'h00000230, 32'h00004820, 32'h000001c0, 32'h00000070, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#281 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h00000230, 32'hxxxxxxxx, 32'h00000070};
#282 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h01254820, 32'h00000244, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000230, 32'h00000014, 32'h00000244, 5'h09, 32'h00000244, 32'h00004820, 32'h00000230, 32'h00000014, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#282 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h00000244, 32'hxxxxxxxx, 32'h00000014};
#283 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h00094880, 32'h00000910, 1'b0, 32'hxxxxxxxx, 32'h00000244, 32'h00000000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000244, 32'h00000910, 5'h09, 32'h00000910, 32'h00004880, 32'h00000002, 32'h00000244, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#283 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h00000910, 32'hxxxxxxxx, 32'h00000244};
#284 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h01094020, 32'h10020910, 1'b0, 32'h00000003, 32'h00000910, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000910, 32'h10020910, 5'h08, 32'h10020910, 32'h00004020, 32'h10020000, 32'h00000910, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#284 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h10020910, 32'h00000003, 32'h00000910};
#284 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h047, 10'h000, 12'hf20};
#284 bmem_addr <= 'h0007;
#285 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'had040000, 32'h10020910, 1'b1, 32'h00000003, 32'h00000002, 32'h00000000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10020910, 32'h00000002, 32'h10020910, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020910, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#285 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h10020910, 32'h00000003, 32'h00000002};
#285 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h047, 10'h000, 12'hf20};
#286 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001d, 32'h008c008c, 32'h10010ffc, 32'h00400024, 32'h00400024};
#286 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h00400024, 32'h00400024, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'h1f, 32'h00400024, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#286 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h047, 10'h000, 12'hf20};
#287 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h10020910, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020910, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#287 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h008c008c, 32'h10010ff8, 32'hxxxxxxxx, 32'h10020910};
#288 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h00000910, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000910, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#288 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h008c008c, 32'h10010ff4, 32'hxxxxxxxx, 32'h00000910};
#288 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h048, 10'h000, 12'hf20};
#288 bmem_addr <= 'h0008;
#289 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000070, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000070, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#289 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h008c008c, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000070};
#290 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#290 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h10011000, 32'h00000000, 32'h10010ff0};
#291 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400144, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0004, 1'b0, 5'bxxxxx, 1'bx, 32'h00400024, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#291 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h008c008c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#292 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h049, 10'h000, 12'hf20};
#292 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h0c1000d3, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0004, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400028, 32'h000000d3, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#292 bmem_addr <= 'h0009;
#292 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h008c008c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#293 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040034c, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001d, 32'h10020000, 32'h00000000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#293 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h10030000, 32'h0000001d, 32'h10020000};
#294 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400350, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001d, 32'h00000000, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#294 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h10030000, 32'h0000001d, 32'h00000000};
#295 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400354, 32'h8c220004, 32'h10030004, 1'b0, 32'h008c008c, 32'h00000003, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000003, 32'h10030004, 5'h02, 32'h008c008c, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#295 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001d, 32'h008c008c, 32'h10030004, 32'h008c008c, 32'h00000003};
#296 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400358, 32'h00021402, 32'h0000008c, 1'b0, 32'hxxxxxxxx, 32'h008c008c, 32'h00000000, 16'h0004, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h008c008c, 32'h0000008c, 5'h02, 32'h0000008c, 32'h00001402, 32'h00000010, 32'h008c008c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#296 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h0000008c, 32'hxxxxxxxx, 32'h008c008c};
#296 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h04a, 10'h000, 12'hf20};
#296 bmem_addr <= 'h000a;
#297 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040035c, 32'h304201ff, 32'h0000008c, 1'b0, 32'hxxxxxxxx, 32'h0000008c, 32'h00000000, 16'h0004, 1'b1, 5'bx0000, 1'b0, 32'h0000008c, 32'h0000008c, 32'h0000008c, 5'h02, 32'h0000008c, 32'h000001ff, 32'h0000008c, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#297 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h0000008c, 32'hxxxxxxxx, 32'h0000008c};
#298 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400360, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0004, 1'b0, 5'bxxxxx, 1'bx, 32'h00400028, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#298 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h008c008c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#299 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h00022300, 32'h0008c000, 1'b0, 32'hxxxxxxxx, 32'h0000008c, 32'h00000000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000008c, 32'h0008c000, 5'h04, 32'h0008c000, 32'h00002300, 32'h0000000c, 32'h0000008c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#299 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h008c008c, 32'h0008c000, 32'hxxxxxxxx, 32'h0000008c};
#300 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00960096, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#300 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h04b, 10'h000, 12'hf20};
#300 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h0c1000de, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0004, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400030, 32'h000000de, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#300 bmem_addr <= 'h000b;
#301 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400378, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001d, 32'h10030000, 32'h00000000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#301 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00960096, 32'h10030000, 32'h0000001d, 32'h10030000};
#302 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040037c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001d, 32'h00000000, 32'h00000000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#302 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00960096, 32'h10030000, 32'h0000001d, 32'h00000000};
#303 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400380, 32'hac240008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h0008c000, 32'h00000000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h0008c000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#303 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001d, 32'h00960096, 32'h10030008, 32'hxxxxxxxx, 32'h0008c000};
#304 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400384, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0008c000, 16'h0004, 1'b0, 5'bxxxxx, 1'bx, 32'h00400030, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#304 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h04c, 10'h000, 12'hf20};
#304 bmem_addr <= 'h000c;
#304 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00960096, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#305 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h0c1000d9, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h0008c000, 16'h0004, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400034, 32'h000000d9, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#305 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00960096, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#306 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400364, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001d, 32'h10030000, 32'h0008c000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#306 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00960096, 32'h10030000, 32'h0000001d, 32'h10030000};
#307 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400368, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001d, 32'h00000000, 32'h0008c000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#307 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00960096, 32'h10030000, 32'h0000001d, 32'h00000000};
#308 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h04d, 10'h000, 12'hf20};
#308 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040036c, 32'h8c220004, 32'h10030004, 1'b0, 32'h00960096, 32'h0000008c, 32'h0008c000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h0000008c, 32'h10030004, 5'h02, 32'h00960096, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#308 bmem_addr <= 'h000d;
#308 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001d, 32'h00960096, 32'h10030004, 32'h00960096, 32'h0000008c};
#309 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400370, 32'h304201ff, 32'h00000096, 1'b0, 32'hxxxxxxxx, 32'h00960096, 32'h0008c000, 16'h0004, 1'b1, 5'bx0000, 1'b0, 32'h00960096, 32'h00960096, 32'h00000096, 5'h02, 32'h00000096, 32'h000001ff, 32'h00960096, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#309 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h0000001d, 32'h00960096, 32'h00000096, 32'hxxxxxxxx, 32'h00960096};
#310 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400374, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0008c000, 16'h0004, 1'b0, 5'bxxxxx, 1'bx, 32'h00400034, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#310 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00960096, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#311 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h00021142, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000096, 32'h0008c000, 16'h0004, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00000096, 32'h00000004, 5'h02, 32'h00000004, 32'h00001142, 32'h00000005, 32'h00000096, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#311 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001d, 32'h00960096, 32'h00000004, 32'hxxxxxxxx, 32'h00000096};
#312 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h24040001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h0008c000, 32'h0008c000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0008c000, 32'h00000001, 5'h04, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#312 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00960096, 32'h00000001, 32'hxxxxxxxx, 32'h0008c000};
#312 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h04e, 10'h000, 12'hf20};
#312 bmem_addr <= 'h000e;
#313 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h00442004, 32'h00000010, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h0008c000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000004, 32'h00000001, 32'h00000010, 5'h04, 32'h00000010, 32'h00002004, 32'h00000004, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#313 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001d, 32'h00960096, 32'h00000010, 32'hxxxxxxxx, 32'h00000001};
#314 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h0c1000e6, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h0008c000, 16'h0004, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400044, 32'h000000e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#314 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00960096, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#315 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400398, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001d, 32'h10030000, 32'h0008c000, 16'h0004, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#315 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00960096, 32'h10030000, 32'h0000001d, 32'h10030000};
#316 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h04f, 10'h000, 12'hf20};
#316 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040039c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001d, 32'h00000000, 32'h0008c000, 16'h0004, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#316 bmem_addr <= 'h000f;
#316 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00960096, 32'h10030000, 32'h0000001d, 32'h00000000};
#317 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a0, 32'hac24000c, 32'h1003000c, 1'b1, 32'hxxxxxxxx, 32'h00000010, 32'h0008c000, 16'h0004, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000010, 32'h1003000c, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10030000, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#317 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b1, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h00960096, 32'h1003000c, 32'hxxxxxxxx, 32'h00000010};
#318 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a4, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0008c000, 16'h0010, 1'b0, 5'bxxxxx, 1'bx, 32'h00400044, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#318 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00960096, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#319 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h2404000f, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000010, 32'h0000000f, 5'h04, 32'h0000000f, 32'h0000000f, 32'h00000000, 32'h0000000f, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#319 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h00960096, 32'h0000000f, 32'hxxxxxxxx, 32'h00000010};
#320 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00a000a0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#320 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h0c100066, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h0008c000, 16'h0010, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h0040004c, 32'h00000066, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#320 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h050, 10'h000, 12'hf20};
#320 smem_addr <= 'h005;
#320 bmem_addr <= 'h0000;
#321 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#321 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00a000a0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#322 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h00400024, 32'h0040004c, 32'h0008c000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#322 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001d, 32'h00a000a0, 32'h10010ffc, 32'h00400024, 32'h0040004c};
#322 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h050, 10'h000, 12'hf20};
#323 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00a000a0, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#323 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0008c000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#324 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h051, 10'h000, 12'hf20};
#324 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0008c000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#324 bmem_addr <= 'h0001;
#324 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00a000a0, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#325 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0008c000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#325 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00a000a0, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#326 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001d, 32'h10030000, 32'h0008c000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#326 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00a000a0, 32'h10030000, 32'h0000001d, 32'h10030000};
#326 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h051, 10'h000, 12'hf20};
#327 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001d, 32'h00000000, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#327 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00a000a0, 32'h10030000, 32'h0000001d, 32'h00000000};
#328 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h052, 10'h000, 12'hf20};
#328 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8c220000, 32'h10030000, 1'b0, 32'h0000001d, 32'h00000004, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000004, 32'h10030000, 5'h02, 32'h0000001d, 32'h00000000, 32'h10030000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#328 bmem_addr <= 'h0002;
#328 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00a000a0, 32'h10030000, 32'h0000001d, 32'h00000004};
#329 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h1040000f, 32'h0000001d, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0008c000, 16'h0010, 1'b0, 5'b1xx01, 1'b0, 32'h0000001d, 32'h00000000, 32'h0000001d, 5'hxx, 32'hxxxxxxxx, 32'h0000000f, 32'h0000001d, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#329 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000004b, 32'h0000001d, 32'h00a000a0, 32'h0000001d, 32'hxxxxxxxx, 32'h00000000};
#330 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h00024821, 32'h0000001d, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001d, 5'h09, 32'h0000001d, 32'h00004821, 32'h00000000, 32'h0000001d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#330 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000004b, 32'h0000001d, 32'h00a000a0, 32'h0000001d, 32'hxxxxxxxx, 32'h0000001d};
#331 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c0, 32'h24020000, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h0000001d, 32'h00000000, 5'h02, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#331 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00a000a0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d};
#332 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c4, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10030000, 32'h0008c000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#332 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00a000a0, 32'h10010000, 32'h00000000, 32'h10030000};
#332 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h053, 10'h000, 12'hf20};
#332 bmem_addr <= 'h0003;
#333 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c8, 32'h34280008, 32'h10010008, 1'b0, 32'h0000001c, 32'hxxxxxxxx, 32'h0008c000, 16'h0010, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010008, 5'h08, 32'h10010008, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#333 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001d, 32'h00a000a0, 32'h10010008, 32'h0000001c, 32'hxxxxxxxx};
#334 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001cc, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h0008c000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#334 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00a000a0, 32'h10010000, 32'h00000000, 32'h10010000};
#335 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d0, 32'h342a0018, 32'h10010018, 1'b0, 32'h0000003b, 32'hxxxxxxxx, 32'h0008c000, 16'h0010, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010018, 5'h0a, 32'h10010018, 32'h00000018, 32'h10010000, 32'h00000018, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#335 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h0000001d, 32'h00a000a0, 32'h10010018, 32'h0000003b, 32'hxxxxxxxx};
#336 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d4, 32'h01485022, 32'h00000010, 1'b0, 32'hxxxxxxxx, 32'h10010008, 32'h0008c000, 16'h0010, 1'b1, 5'b1xx01, 1'b0, 32'h10010018, 32'h10010008, 32'h00000010, 5'h0a, 32'h00000010, 32'h00005022, 32'h10010018, 32'h10010008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#336 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001d, 32'h00a000a0, 32'h00000010, 32'hxxxxxxxx, 32'h10010008};
#336 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h054, 10'h000, 12'hf20};
#336 bmem_addr <= 'h0004;
#337 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h0008c000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#337 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00a000a0, 32'h10010000, 32'h00000000, 32'h10010000};
#338 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#338 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00a000a0, 32'h10010000, 32'h00000000, 32'h00000000};
#339 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010008, 1'b0, 32'h0000001c, 32'h10010008, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h10010008, 32'h10010008, 5'h08, 32'h0000001c, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#339 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001d, 32'h00a000a0, 32'h10010008, 32'h0000001c, 32'h10010008};
#340 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001d, 32'h00aa00aa, 32'h00000004, 32'hxxxxxxxx, 32'h00000000};
#340 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000004, 5'h02, 32'h00000004, 32'h00000004, 32'h00000000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#340 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h055, 10'h000, 12'hf20};
#340 bmem_addr <= 'h0005;
#341 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'hffffffff, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0008c000, 16'h0010, 1'b0, 5'b1xx01, 1'b0, 32'h0000001c, 32'h0000001d, 32'hffffffff, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001c, 32'h0000001d, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#341 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001d, 32'h00aa00aa, 32'hffffffff, 32'hxxxxxxxx, 32'h0000001d};
#342 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0008c000, 16'h0010, 1'b1, 5'b1x011, 1'b0, 32'h00000004, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h00000004, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#342 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00aa00aa, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#343 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0008c000, 16'h0010, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#343 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00aa00aa, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#344 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h056, 10'h000, 12'hf20};
#344 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h0008c000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#344 bmem_addr <= 'h0006;
#344 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00aa00aa, 32'h10010000, 32'h00000000, 32'h00000001};
#345 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010004, 1'b0, 32'h00000003, 32'h00000004, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000004, 32'h10010004, 5'h01, 32'h10010004, 32'h00000821, 32'h10010000, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#345 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001d, 32'h00aa00aa, 32'h10010004, 32'h00000003, 32'h00000004};
#346 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h1001000c, 1'b0, 32'h00000023, 32'h0000001c, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010004, 32'h0000001c, 32'h1001000c, 5'h08, 32'h00000023, 32'h00000008, 32'h10010004, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#346 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h00aa00aa, 32'h1001000c, 32'h00000023, 32'h0000001c};
#347 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000008, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000004, 32'h00000004, 32'h00000008, 5'h02, 32'h00000008, 32'h00000004, 32'h00000004, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#347 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001d, 32'h00aa00aa, 32'h00000008, 32'hxxxxxxxx, 32'h00000004};
#348 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000006, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0008c000, 16'h0010, 1'b0, 5'b1xx01, 1'b0, 32'h00000023, 32'h0000001d, 32'h00000006, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h00000023, 32'h0000001d, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#348 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001d, 32'h00aa00aa, 32'h00000006, 32'hxxxxxxxx, 32'h0000001d};
#348 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h057, 10'h000, 12'hf20};
#348 bmem_addr <= 'h0007;
#349 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0008c000, 16'h0010, 1'b1, 5'b1x011, 1'b0, 32'h00000008, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h00000008, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#349 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00aa00aa, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#350 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0008c000, 16'h0010, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#350 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00aa00aa, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#351 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h0008c000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#351 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00aa00aa, 32'h10010000, 32'h00000000, 32'h00000001};
#352 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010008, 1'b0, 32'h0000001c, 32'h00000008, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000008, 32'h10010008, 5'h01, 32'h10010008, 32'h00000821, 32'h10010000, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#352 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001d, 32'h00aa00aa, 32'h10010008, 32'h0000001c, 32'h00000008};
#352 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h058, 10'h000, 12'hf20};
#352 bmem_addr <= 'h0008;
#353 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010010, 1'b0, 32'h0000001d, 32'h00000023, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010008, 32'h00000023, 32'h10010010, 5'h08, 32'h0000001d, 32'h00000008, 32'h10010008, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#353 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001d, 32'h00aa00aa, 32'h10010010, 32'h0000001d, 32'h00000023};
#354 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h0000000c, 1'b0, 32'hxxxxxxxx, 32'h00000008, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000008, 32'h00000008, 32'h0000000c, 5'h02, 32'h0000000c, 32'h00000004, 32'h00000008, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#354 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h00aa00aa, 32'h0000000c, 32'hxxxxxxxx, 32'h00000008};
#355 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0008c000, 16'h0010, 1'b0, 5'b1xx01, 1'b1, 32'h0000001d, 32'h0000001d, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001d, 32'h0000001d, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#355 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00aa00aa, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d};
#356 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h059, 10'h000, 12'hf20};
#356 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f8, 32'h00021082, 32'h00000003, 1'b0, 32'hxxxxxxxx, 32'h0000000c, 32'h0008c000, 16'h0010, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h0000000c, 32'h00000003, 5'h02, 32'h00000003, 32'h00001082, 32'h00000002, 32'h0000000c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#356 bmem_addr <= 'h0009;
#356 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00aa00aa, 32'h00000003, 32'hxxxxxxxx, 32'h0000000c};
#357 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001fc, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h0040004c, 32'h0040004c, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'h1f, 32'h0040004c, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#357 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h0000001d, 32'h00aa00aa, 32'h10010ffc, 32'h0040004c, 32'h0040004c};
#358 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400200, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001d, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#358 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00aa00aa, 32'h10010ff8, 32'hxxxxxxxx, 32'h0000001d};
#359 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400204, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h0000001d, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001d, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#359 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00aa00aa, 32'h10010ff4, 32'hxxxxxxxx, 32'h0000001d};
#360 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00b400b4, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000010};
#360 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400208, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000010, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#360 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h05a, 10'h000, 12'hf20};
#360 bmem_addr <= 'h000a;
#361 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040020c, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#361 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00b400b4, 32'h10011000, 32'h00000000, 32'h10010ff0};
#362 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400210, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0008c000, 16'h0010, 1'b0, 5'bxxxxx, 1'bx, 32'h0040004c, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#362 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00b400b4, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#363 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h00028021, 32'h00000003, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000003, 5'h10, 32'h00000003, 32'hxxxx8021, 32'h00000000, 32'h00000003, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#363 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00b400b4, 32'h00000003, 32'hxxxxxxxx, 32'h00000003};
#364 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h05b, 10'h000, 12'hf20};
#364 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h0c1000e2, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h0008c000, 16'h0010, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400054, 32'h000000e2, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#364 bmem_addr <= 'h000b;
#364 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00b400b4, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#365 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400388, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001d, 32'h10010008, 32'h0008c000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010008, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#365 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00b400b4, 32'h10030000, 32'h0000001d, 32'h10010008};
#366 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040038c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001d, 32'h00000000, 32'h0008c000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#366 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00b400b4, 32'h10030000, 32'h0000001d, 32'h00000000};
#367 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400390, 32'hac200008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h00000000, 32'h0008c000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#367 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001d, 32'h00b400b4, 32'h10030008, 32'hxxxxxxxx, 32'h00000000};
#368 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400394, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0010, 1'b0, 5'bxxxxx, 1'bx, 32'h00400054, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#368 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h05c, 10'h000, 12'hf20};
#368 bmem_addr <= 'h000c;
#368 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00b400b4, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#369 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400054, 32'h1200ffef, 32'h00000003, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0010, 1'b0, 5'b1xx01, 1'b0, 32'h00000003, 32'h00000000, 32'h00000003, 5'hxx, 32'hxxxxxxxx, 32'hffffffef, 32'h00000003, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#369 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00b400b4, 32'h00000003, 32'hxxxxxxxx, 32'h00000000};
#370 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400058, 32'h20010001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h10030000, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h10030000, 32'h00000001, 5'h01, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#370 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00b400b4, 32'h00000001, 32'hxxxxxxxx, 32'h10030000};
#371 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040005c, 32'h14300005, 32'hfffffffe, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0010, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000003, 32'hfffffffe, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000001, 32'h00000003, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#371 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001d, 32'h00b400b4, 32'hfffffffe, 32'hxxxxxxxx, 32'h00000003};
#372 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h05d, 10'h000, 12'hf20};
#372 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400074, 32'h20010002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000001, 32'h00000002, 5'h01, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#372 bmem_addr <= 'h000d;
#372 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00b400b4, 32'h00000002, 32'hxxxxxxxx, 32'h00000001};
#373 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400078, 32'h14300005, 32'hffffffff, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0010, 1'b0, 5'b1xx01, 1'b0, 32'h00000002, 32'h00000003, 32'hffffffff, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000002, 32'h00000003, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#373 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001d, 32'h00b400b4, 32'hffffffff, 32'hxxxxxxxx, 32'h00000003};
#374 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400090, 32'h20010003, 32'h00000003, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000003, 5'h01, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#374 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00b400b4, 32'h00000003, 32'hxxxxxxxx, 32'h00000002};
#375 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400094, 32'h14300005, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0010, 1'b0, 5'b1xx01, 1'b1, 32'h00000003, 32'h00000003, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000003, 32'h00000003, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#375 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00b400b4, 32'h00000000, 32'hxxxxxxxx, 32'h00000003};
#376 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h05e, 10'h000, 12'hf20};
#376 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400098, 32'h2252ffff, 32'h0000000d, 1'b0, 32'hxxxxxxxx, 32'h0000000e, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h0000000e, 32'h0000000e, 32'h0000000d, 5'h12, 32'h0000000d, 32'hffffffff, 32'h0000000e, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#376 bmem_addr <= 'h000e;
#376 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h00b400b4, 32'h0000000d, 32'hxxxxxxxx, 32'h0000000e};
#377 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040009c, 32'h0240082a, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0010, 1'b1, 5'b1x011, 1'b1, 32'h0000000d, 32'h00000000, 32'h00000000, 5'h01, 32'h00000000, 32'h0000082a, 32'h0000000d, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#377 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00b400b4, 32'h00000000, 32'hxxxxxxxx, 32'h00000000};
#378 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000a0, 32'h1020ffdc, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0010, 1'b0, 5'b1xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'hffffffdc, 32'h00000000, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#379 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h24040002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#379 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00b400b4, 32'h00000002, 32'hxxxxxxxx, 32'h0000000f};
#380 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h0000001d, 32'h00be00be, 32'h00000014, 32'hxxxxxxxx, 32'h00000014};
#380 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00112821, 32'h00000014, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000014, 32'h00000014, 5'h05, 32'h00000014, 32'h00002821, 32'h00000000, 32'h00000014, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#380 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h05f, 10'h000, 12'hf20};
#380 bmem_addr <= 'h000f;
#381 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h00123021, 32'h0000000d, 1'b0, 32'hxxxxxxxx, 32'h0000000d, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000d, 32'h0000000d, 5'h06, 32'h0000000d, 32'h00003021, 32'h00000000, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#381 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001d, 32'h00be00be, 32'h0000000d, 32'hxxxxxxxx, 32'h0000000d};
#382 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h0c10003e, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0010, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400024, 32'h0000003e, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#382 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001d, 32'h00be00be, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#383 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000f8, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#383 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00be00be, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#384 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h0040004c, 32'h00400024, 32'h00000000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#384 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h0000001d, 32'h00be00be, 32'h10010ffc, 32'h0040004c, 32'h00400024};
#384 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h060, 10'h000, 12'h0f0};
#384 smem_addr <= 'h006;
#384 bmem_addr <= 'h0100;
#384 charcode  <= 'h01;
#385 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00be00be, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#385 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#386 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#386 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00be00be, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#387 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#387 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00be00be, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#388 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h061, 10'h000, 12'h0f0};
#388 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#388 bmem_addr <= 'h0101;
#388 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00be00be, 32'h10020000, 32'h00000000, 32'h00000000};
#389 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0010, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'hxxxxxxxx, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#389 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00be00be, 32'h10020000, 32'h00000000, 32'hxxxxxxxx};
#390 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h00064940, 32'h000001a0, 1'b0, 32'hxxxxxxxx, 32'h0000000d, 32'h00000000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000d, 32'h000001a0, 5'h09, 32'h000001a0, 32'h00004940, 32'h00000005, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#390 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00be00be, 32'h000001a0, 32'hxxxxxxxx, 32'h0000000d};
#391 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h000650c0, 32'h00000068, 1'b0, 32'hxxxxxxxx, 32'h0000000d, 32'h00000000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000068, 5'h0a, 32'h00000068, 32'h000050c0, 32'h00000003, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#391 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h0000001d, 32'h00be00be, 32'h00000068, 32'hxxxxxxxx, 32'h0000000d};
#392 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h062, 10'h000, 12'h0f0};
#392 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h012a4820, 32'h00000208, 1'b0, 32'hxxxxxxxx, 32'h00000068, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h000001a0, 32'h00000068, 32'h00000208, 5'h09, 32'h00000208, 32'h00004820, 32'h000001a0, 32'h00000068, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#392 bmem_addr <= 'h0102;
#392 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h0000001d, 32'h00be00be, 32'h00000208, 32'hxxxxxxxx, 32'h00000068};
#393 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h01254820, 32'h0000021c, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000208, 32'h00000014, 32'h0000021c, 5'h09, 32'h0000021c, 32'h00004820, 32'h00000208, 32'h00000014, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#393 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h0000001d, 32'h00be00be, 32'h0000021c, 32'hxxxxxxxx, 32'h00000014};
#394 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h00094880, 32'h00000870, 1'b0, 32'hxxxxxxxx, 32'h0000021c, 32'h00000000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000021c, 32'h00000870, 5'h09, 32'h00000870, 32'h00004880, 32'h00000002, 32'h0000021c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#394 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00be00be, 32'h00000870, 32'hxxxxxxxx, 32'h0000021c};
#395 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h01094020, 32'h10020870, 1'b0, 32'h00000000, 32'h00000870, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000870, 32'h10020870, 5'h08, 32'h10020870, 32'h00004020, 32'h10020000, 32'h00000870, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#395 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00be00be, 32'h10020870, 32'h00000000, 32'h00000870};
#396 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'had040000, 32'h10020870, 1'b1, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10020870, 32'h00000002, 32'h10020870, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020870, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#396 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001d, 32'h00be00be, 32'h10020870, 32'h00000000, 32'h00000002};
#396 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h063, 10'h000, 12'h0f0};
#396 bmem_addr <= 'h0103;
#397 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001d, 32'h00be00be, 32'h10010ffc, 32'h00400024, 32'h00400024};
#397 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h00400024, 32'h00400024, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'h1f, 32'h00400024, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#397 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h063, 10'h000, 12'h0f0};
#398 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h10020870, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020870, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#398 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00be00be, 32'h10010ff8, 32'hxxxxxxxx, 32'h10020870};
#399 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h00000870, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000870, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#399 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001d, 32'h00be00be, 32'h10010ff4, 32'hxxxxxxxx, 32'h00000870};
#400 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00c800c8, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000068};
#400 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000068, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000068, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#400 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h064, 10'h000, 12'h0f0};
#400 bmem_addr <= 'h0104;
#401 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#401 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00c800c8, 32'h10011000, 32'h00000000, 32'h10010ff0};
#402 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400144, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0010, 1'b0, 5'bxxxxx, 1'bx, 32'h00400024, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#402 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00c800c8, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#403 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h0c1000d3, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0010, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400028, 32'h000000d3, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#403 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00c800c8, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#404 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040034c, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10020000, 32'h00000000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#404 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h065, 10'h000, 12'h0f0};
#404 bmem_addr <= 'h0105;
#404 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00c800c8, 32'h10030000, 32'h00000023, 32'h10020000};
#405 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400350, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#405 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00c800c8, 32'h10030000, 32'h00000023, 32'h00000000};
#406 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400354, 32'h8c220004, 32'h10030004, 1'b0, 32'h00c800c8, 32'h00000003, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000003, 32'h10030004, 5'h02, 32'h00c800c8, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#406 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000023, 32'h00c800c8, 32'h10030004, 32'h00c800c8, 32'h00000003};
#407 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400358, 32'h00021402, 32'h000000c8, 1'b0, 32'hxxxxxxxx, 32'h00c800c8, 32'h00000000, 16'h0010, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00c800c8, 32'h000000c8, 5'h02, 32'h000000c8, 32'h00001402, 32'h00000010, 32'h00c800c8, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#407 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00c800c8, 32'h000000c8, 32'hxxxxxxxx, 32'h00c800c8};
#408 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040035c, 32'h304201ff, 32'h000000c8, 1'b0, 32'hxxxxxxxx, 32'h000000c8, 32'h00000000, 16'h0010, 1'b1, 5'bx0000, 1'b0, 32'h000000c8, 32'h000000c8, 32'h000000c8, 5'h02, 32'h000000c8, 32'h000001ff, 32'h000000c8, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#408 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00c800c8, 32'h000000c8, 32'hxxxxxxxx, 32'h000000c8};
#408 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h066, 10'h000, 12'h0f0};
#408 bmem_addr <= 'h0106;
#409 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400360, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0010, 1'b0, 5'bxxxxx, 1'bx, 32'h00400028, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#409 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00c800c8, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#410 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h00022300, 32'h000c8000, 1'b0, 32'hxxxxxxxx, 32'h000000c8, 32'h00000000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000000c8, 32'h000c8000, 5'h04, 32'h000c8000, 32'h00002300, 32'h0000000c, 32'h000000c8, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#410 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00c800c8, 32'h000c8000, 32'hxxxxxxxx, 32'h000000c8};
#411 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h0c1000de, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0010, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400030, 32'h000000de, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#411 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00c800c8, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#412 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400378, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10030000, 32'h00000000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#412 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h067, 10'h000, 12'h0f0};
#412 bmem_addr <= 'h0107;
#412 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00c800c8, 32'h10030000, 32'h00000023, 32'h10030000};
#413 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040037c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h00000000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#413 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00c800c8, 32'h10030000, 32'h00000023, 32'h00000000};
#414 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400380, 32'hac240008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h000c8000, 32'h00000000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h000c8000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#414 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000023, 32'h00c800c8, 32'h10030008, 32'hxxxxxxxx, 32'h000c8000};
#415 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400384, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000c8000, 16'h0010, 1'b0, 5'bxxxxx, 1'bx, 32'h00400030, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#415 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00c800c8, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#416 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h068, 10'h000, 12'h0f0};
#416 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h0c1000d9, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h000c8000, 16'h0010, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400034, 32'h000000d9, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#416 bmem_addr <= 'h0108;
#416 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00c800c8, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#417 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400364, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10030000, 32'h000c8000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#417 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00c800c8, 32'h10030000, 32'h00000023, 32'h10030000};
#418 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400368, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h000c8000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#418 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00c800c8, 32'h10030000, 32'h00000023, 32'h00000000};
#419 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040036c, 32'h8c220004, 32'h10030004, 1'b0, 32'h00c800c8, 32'h000000c8, 32'h000c8000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h000000c8, 32'h10030004, 5'h02, 32'h00c800c8, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#419 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000023, 32'h00c800c8, 32'h10030004, 32'h00c800c8, 32'h000000c8};
#420 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00d200d2, 32'h000000d2, 32'hxxxxxxxx, 32'h00d200d2};
#420 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400370, 32'h304201ff, 32'h000000d2, 1'b0, 32'hxxxxxxxx, 32'h00d200d2, 32'h000c8000, 16'h0010, 1'b1, 5'bx0000, 1'b0, 32'h00d200d2, 32'h00d200d2, 32'h000000d2, 5'h02, 32'h000000d2, 32'h000001ff, 32'h00d200d2, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#420 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h069, 10'h000, 12'h0f0};
#420 bmem_addr <= 'h0109;
#421 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400374, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000c8000, 16'h0010, 1'b0, 5'bxxxxx, 1'bx, 32'h00400034, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#421 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00d200d2, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#422 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h00021142, 32'h00000006, 1'b0, 32'hxxxxxxxx, 32'h000000d2, 32'h000c8000, 16'h0010, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h000000d2, 32'h00000006, 5'h02, 32'h00000006, 32'h00001142, 32'h00000005, 32'h000000d2, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#422 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000023, 32'h00d200d2, 32'h00000006, 32'hxxxxxxxx, 32'h000000d2};
#423 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h24040001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h000c8000, 32'h000c8000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h000c8000, 32'h00000001, 5'h04, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#423 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00d200d2, 32'h00000001, 32'hxxxxxxxx, 32'h000c8000};
#424 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h00442004, 32'h00000040, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h000c8000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000006, 32'h00000001, 32'h00000040, 5'h04, 32'h00000040, 32'h00002004, 32'h00000006, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#424 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h00000023, 32'h00d200d2, 32'h00000040, 32'hxxxxxxxx, 32'h00000001};
#424 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h06a, 10'h000, 12'h0f0};
#424 bmem_addr <= 'h010a;
#425 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h0c1000e6, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h000c8000, 16'h0010, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h00400044, 32'h000000e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#425 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00d200d2, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#426 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400398, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10030000, 32'h000c8000, 16'h0010, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#426 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00d200d2, 32'h10030000, 32'h00000023, 32'h10030000};
#427 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040039c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h000c8000, 16'h0010, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#427 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00d200d2, 32'h10030000, 32'h00000023, 32'h00000000};
#428 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h06b, 10'h000, 12'h0f0};
#428 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a0, 32'hac24000c, 32'h1003000c, 1'b1, 32'hxxxxxxxx, 32'h00000040, 32'h000c8000, 16'h0010, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000040, 32'h1003000c, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10030000, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#428 bmem_addr <= 'h010b;
#428 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b1, 32'h00000003, 32'h00000023, 32'h00000023, 32'h00d200d2, 32'h1003000c, 32'hxxxxxxxx, 32'h00000040};
#429 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a4, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000c8000, 16'h0040, 1'b0, 5'bxxxxx, 1'bx, 32'h00400044, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#429 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00d200d2, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#430 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h2404000f, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h00000040, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000040, 32'h0000000f, 5'h04, 32'h0000000f, 32'h0000000f, 32'h00000000, 32'h0000000f, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#430 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000023, 32'h00d200d2, 32'h0000000f, 32'hxxxxxxxx, 32'h00000040};
#431 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h0c100066, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h000c8000, 16'h0040, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000003, 32'hxxxxxxxx, 5'h1f, 32'h0040004c, 32'h00000066, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#431 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00d200d2, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000003};
#432 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#432 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h06c, 10'h000, 12'h0f0};
#432 bmem_addr <= 'h010c;
#432 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00d200d2, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#433 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h00400024, 32'h0040004c, 32'h000c8000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#433 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h00000023, 32'h00d200d2, 32'h10010ffc, 32'h00400024, 32'h0040004c};
#433 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h06c, 10'h000, 12'h0f0};
#434 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00d200d2, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#434 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h000c8000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#435 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h000c8000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#435 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00d200d2, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#436 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h06d, 10'h000, 12'h0f0};
#436 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h000c8000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#436 bmem_addr <= 'h010d;
#436 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00d200d2, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#437 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10030000, 32'h000c8000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#437 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00d200d2, 32'h10030000, 32'h00000023, 32'h10030000};
#437 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h06d, 10'h000, 12'h0f0};
#438 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#438 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00d200d2, 32'h10030000, 32'h00000023, 32'h00000000};
#439 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8c220000, 32'h10030000, 1'b0, 32'h00000023, 32'h00000006, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000006, 32'h10030000, 5'h02, 32'h00000023, 32'h00000000, 32'h10030000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#439 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00d200d2, 32'h10030000, 32'h00000023, 32'h00000006};
#440 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000043, 32'h00000023, 32'h00dc00dc, 32'h00000023, 32'hxxxxxxxx, 32'h00000000};
#440 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h1040000f, 32'h00000023, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000c8000, 16'h0040, 1'b0, 5'b1xx01, 1'b0, 32'h00000023, 32'h00000000, 32'h00000023, 5'hxx, 32'hxxxxxxxx, 32'h0000000f, 32'h00000023, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#440 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h06e, 10'h000, 12'h0f0};
#440 bmem_addr <= 'h010e;
#441 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h00024821, 32'h00000023, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000023, 32'h00000023, 5'h09, 32'h00000023, 32'h00004821, 32'h00000000, 32'h00000023, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#441 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000043, 32'h00000023, 32'h00dc00dc, 32'h00000023, 32'hxxxxxxxx, 32'h00000023};
#442 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c0, 32'h24020000, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000023, 32'h00000000, 5'h02, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#442 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00dc00dc, 32'h00000000, 32'hxxxxxxxx, 32'h00000023};
#443 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c4, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10030000, 32'h000c8000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#443 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00dc00dc, 32'h10010000, 32'h00000000, 32'h10030000};
#444 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c8, 32'h34280008, 32'h10010008, 1'b0, 32'h0000001c, 32'hxxxxxxxx, 32'h000c8000, 16'h0040, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010008, 5'h08, 32'h10010008, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#444 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000023, 32'h00dc00dc, 32'h10010008, 32'h0000001c, 32'hxxxxxxxx};
#444 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h06f, 10'h000, 12'h0f0};
#444 bmem_addr <= 'h010f;
#445 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001cc, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h000c8000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#445 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00dc00dc, 32'h10010000, 32'h00000000, 32'h10010000};
#446 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d0, 32'h342a0018, 32'h10010018, 1'b0, 32'h0000003b, 32'hxxxxxxxx, 32'h000c8000, 16'h0040, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010018, 5'h0a, 32'h10010018, 32'h00000018, 32'h10010000, 32'h00000018, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#446 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h00000023, 32'h00dc00dc, 32'h10010018, 32'h0000003b, 32'hxxxxxxxx};
#447 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d4, 32'h01485022, 32'h00000010, 1'b0, 32'hxxxxxxxx, 32'h10010008, 32'h000c8000, 16'h0040, 1'b1, 5'b1xx01, 1'b0, 32'h10010018, 32'h10010008, 32'h00000010, 5'h0a, 32'h00000010, 32'h00005022, 32'h10010018, 32'h10010008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#447 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h00000023, 32'h00dc00dc, 32'h00000010, 32'hxxxxxxxx, 32'h10010008};
#448 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h000c8000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#448 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00dc00dc, 32'h10010000, 32'h00000000, 32'h10010000};
#448 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h070, 10'h000, 12'hfff};
#448 smem_addr <= 'h007;
#448 bmem_addr <= 'h0200;
#448 charcode  <= 'h02;
#449 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#449 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00dc00dc, 32'h10010000, 32'h00000000, 32'h00000000};
#450 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010008, 1'b0, 32'h0000001c, 32'h10010008, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h10010008, 32'h10010008, 5'h08, 32'h0000001c, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#450 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000023, 32'h00dc00dc, 32'h10010008, 32'h0000001c, 32'h10010008};
#451 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000004, 5'h02, 32'h00000004, 32'h00000004, 32'h00000000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#451 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000023, 32'h00dc00dc, 32'h00000004, 32'hxxxxxxxx, 32'h00000000};
#452 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'hfffffff9, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000c8000, 16'h0040, 1'b0, 5'b1xx01, 1'b0, 32'h0000001c, 32'h00000023, 32'hfffffff9, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001c, 32'h00000023, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#452 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00dc00dc, 32'hfffffff9, 32'hxxxxxxxx, 32'h00000023};
#452 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h071, 10'h000, 12'hfff};
#452 bmem_addr <= 'h0201;
#453 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h000c8000, 16'h0040, 1'b1, 5'b1x011, 1'b0, 32'h00000004, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h00000004, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#453 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00dc00dc, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#454 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000c8000, 16'h0040, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#454 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00dc00dc, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#455 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h000c8000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#455 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00dc00dc, 32'h10010000, 32'h00000000, 32'h00000001};
#456 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010004, 1'b0, 32'h00000003, 32'h00000004, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000004, 32'h10010004, 5'h01, 32'h10010004, 32'h00000821, 32'h10010000, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#456 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000023, 32'h00dc00dc, 32'h10010004, 32'h00000003, 32'h00000004};
#456 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h072, 10'h000, 12'hfff};
#456 bmem_addr <= 'h0202;
#457 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h1001000c, 1'b0, 32'h00000023, 32'h0000001c, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010004, 32'h0000001c, 32'h1001000c, 5'h08, 32'h00000023, 32'h00000008, 32'h10010004, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#457 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000023, 32'h00dc00dc, 32'h1001000c, 32'h00000023, 32'h0000001c};
#458 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000008, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000004, 32'h00000004, 32'h00000008, 5'h02, 32'h00000008, 32'h00000004, 32'h00000004, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#458 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000023, 32'h00dc00dc, 32'h00000008, 32'hxxxxxxxx, 32'h00000004};
#459 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000c8000, 16'h0040, 1'b0, 5'b1xx01, 1'b1, 32'h00000023, 32'h00000023, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h00000023, 32'h00000023, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#459 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00dc00dc, 32'h00000000, 32'hxxxxxxxx, 32'h00000023};
#460 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00e600e6, 32'h00000002, 32'hxxxxxxxx, 32'h00000008};
#460 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h073, 10'h000, 12'hfff};
#460 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f8, 32'h00021082, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000008, 32'h000c8000, 16'h0040, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00000008, 32'h00000002, 5'h02, 32'h00000002, 32'h00001082, 32'h00000002, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#460 bmem_addr <= 'h0203;
#461 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001fc, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h0040004c, 32'h0040004c, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'h1f, 32'h0040004c, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#461 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h00000023, 32'h00e600e6, 32'h10010ffc, 32'h0040004c, 32'h0040004c};
#462 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400200, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000023, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#462 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00e600e6, 32'h10010ff8, 32'hxxxxxxxx, 32'h00000023};
#463 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400204, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000023, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#463 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00e600e6, 32'h10010ff4, 32'hxxxxxxxx, 32'h00000023};
#464 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400208, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000010, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#464 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00e600e6, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000010};
#464 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hd, 4'hc, 10'h074, 10'h000, 12'hfdc};
#464 bmem_addr <= 'h0204;
#465 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040020c, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#465 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00e600e6, 32'h10011000, 32'h00000000, 32'h10010ff0};
#466 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400210, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000c8000, 16'h0040, 1'b0, 5'bxxxxx, 1'bx, 32'h0040004c, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#466 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00e600e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#467 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h00028021, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000002, 5'h10, 32'h00000002, 32'hxxxx8021, 32'h00000000, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#467 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00e600e6, 32'h00000002, 32'hxxxxxxxx, 32'h00000002};
#468 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h8, 10'h075, 10'h000, 12'hfc8};
#468 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h0c1000e2, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h000c8000, 16'h0040, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400054, 32'h000000e2, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#468 bmem_addr <= 'h0205;
#468 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00e600e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#469 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400388, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10010004, 32'h000c8000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010004, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#469 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00e600e6, 32'h10030000, 32'h00000023, 32'h10010004};
#470 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040038c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h000c8000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#470 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00e600e6, 32'h10030000, 32'h00000023, 32'h00000000};
#471 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400390, 32'hac200008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h00000000, 32'h000c8000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#471 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000023, 32'h00e600e6, 32'h10030008, 32'hxxxxxxxx, 32'h00000000};
#472 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400394, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0040, 1'b0, 5'bxxxxx, 1'bx, 32'h00400054, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#472 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h076, 10'h000, 12'hfc6};
#472 bmem_addr <= 'h0206;
#472 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00e600e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#473 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400054, 32'h1200ffef, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0040, 1'b0, 5'b1xx01, 1'b0, 32'h00000002, 32'h00000000, 32'h00000002, 5'hxx, 32'hxxxxxxxx, 32'hffffffef, 32'h00000002, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#473 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00e600e6, 32'h00000002, 32'hxxxxxxxx, 32'h00000000};
#474 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400058, 32'h20010001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h10030000, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h10030000, 32'h00000001, 5'h01, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#474 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00e600e6, 32'h00000001, 32'hxxxxxxxx, 32'h10030000};
#475 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040005c, 32'h14300005, 32'hffffffff, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0040, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000002, 32'hffffffff, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000001, 32'h00000002, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#475 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h00000023, 32'h00e600e6, 32'hffffffff, 32'hxxxxxxxx, 32'h00000002};
#476 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h077, 10'h000, 12'hfc6};
#476 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400074, 32'h20010002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000001, 32'h00000002, 5'h01, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#476 bmem_addr <= 'h0207;
#476 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00e600e6, 32'h00000002, 32'hxxxxxxxx, 32'h00000001};
#477 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400078, 32'h14300005, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0040, 1'b0, 5'b1xx01, 1'b1, 32'h00000002, 32'h00000002, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000002, 32'h00000002, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#477 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00e600e6, 32'h00000000, 32'hxxxxxxxx, 32'h00000002};
#478 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040007c, 32'h22310001, 32'h00000015, 1'b0, 32'hxxxxxxxx, 32'h00000014, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000014, 32'h00000014, 32'h00000015, 5'h11, 32'h00000015, 32'h00000001, 32'h00000014, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#478 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h00000023, 32'h00e600e6, 32'h00000015, 32'hxxxxxxxx, 32'h00000014};
#479 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400080, 32'h2a210028, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0040, 1'b1, 5'b1x011, 1'b0, 32'h00000015, 32'h00000002, 32'h00000001, 5'h01, 32'h00000001, 32'h00000028, 32'h00000015, 32'h00000028, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#479 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00e600e6, 32'h00000001, 32'hxxxxxxxx, 32'h00000002};
#480 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00f000f0, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#480 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400084, 32'h1420ffe3, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0040, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hffffffe3, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#480 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h078, 10'h000, 12'hfc6};
#480 bmem_addr <= 'h0208;
#481 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h24040002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#481 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00f000f0, 32'h00000002, 32'hxxxxxxxx, 32'h0000000f};
#482 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00112821, 32'h00000015, 1'b0, 32'hxxxxxxxx, 32'h00000015, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000015, 32'h00000015, 5'h05, 32'h00000015, 32'h00002821, 32'h00000000, 32'h00000015, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#482 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h00000023, 32'h00f000f0, 32'h00000015, 32'hxxxxxxxx, 32'h00000015};
#483 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h00123021, 32'h0000000d, 1'b0, 32'hxxxxxxxx, 32'h0000000d, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000d, 32'h0000000d, 5'h06, 32'h0000000d, 32'h00003021, 32'h00000000, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#483 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000023, 32'h00f000f0, 32'h0000000d, 32'hxxxxxxxx, 32'h0000000d};
#484 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h079, 10'h000, 12'hfc6};
#484 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h0c10003e, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0040, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400024, 32'h0000003e, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#484 bmem_addr <= 'h0209;
#484 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00f000f0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#485 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000f8, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#485 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00f000f0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#486 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h0040004c, 32'h00400024, 32'h00000000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#486 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h00000023, 32'h00f000f0, 32'h10010ffc, 32'h0040004c, 32'h00400024};
#486 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h079, 10'h000, 12'hfc6};
#487 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00f000f0, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#487 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#488 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h8, 10'h07a, 10'h000, 12'hfc8};
#488 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#488 bmem_addr <= 'h020a;
#488 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00f000f0, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#489 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#489 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00f000f0, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#490 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#490 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00f000f0, 32'h10020000, 32'h00000000, 32'h00000001};
#490 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h8, 10'h07a, 10'h000, 12'hfc8};
#491 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0040, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'hxxxxxxxx, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#491 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00f000f0, 32'h10020000, 32'h00000000, 32'hxxxxxxxx};
#492 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h00064940, 32'h000001a0, 1'b0, 32'hxxxxxxxx, 32'h0000000d, 32'h00000000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000d, 32'h000001a0, 5'h09, 32'h000001a0, 32'h00004940, 32'h00000005, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#492 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00f000f0, 32'h000001a0, 32'hxxxxxxxx, 32'h0000000d};
#492 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'he, 4'hc, 10'h07b, 10'h000, 12'hfec};
#492 bmem_addr <= 'h020b;
#493 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h000650c0, 32'h00000068, 1'b0, 32'hxxxxxxxx, 32'h0000000d, 32'h00000000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000068, 5'h0a, 32'h00000068, 32'h000050c0, 32'h00000003, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#493 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h00000023, 32'h00f000f0, 32'h00000068, 32'hxxxxxxxx, 32'h0000000d};
#494 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h012a4820, 32'h00000208, 1'b0, 32'hxxxxxxxx, 32'h00000068, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h000001a0, 32'h00000068, 32'h00000208, 5'h09, 32'h00000208, 32'h00004820, 32'h000001a0, 32'h00000068, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#494 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h00000023, 32'h00f000f0, 32'h00000208, 32'hxxxxxxxx, 32'h00000068};
#495 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h01254820, 32'h0000021d, 1'b0, 32'hxxxxxxxx, 32'h00000015, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000208, 32'h00000015, 32'h0000021d, 5'h09, 32'h0000021d, 32'h00004820, 32'h00000208, 32'h00000015, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#495 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000023, 32'h00f000f0, 32'h0000021d, 32'hxxxxxxxx, 32'h00000015};
#496 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h00094880, 32'h00000874, 1'b0, 32'hxxxxxxxx, 32'h0000021d, 32'h00000000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000021d, 32'h00000874, 5'h09, 32'h00000874, 32'h00004880, 32'h00000002, 32'h0000021d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#496 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000000, 32'h00000023, 32'h00f000f0, 32'h00000874, 32'hxxxxxxxx, 32'h0000021d};
#496 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h07c, 10'h000, 12'hfff};
#496 bmem_addr <= 'h020c;
#497 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h01094020, 32'h10020874, 1'b0, 32'h00000003, 32'h00000874, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000874, 32'h10020874, 5'h08, 32'h10020874, 32'h00004020, 32'h10020000, 32'h00000874, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#497 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000000, 32'h00000023, 32'h00f000f0, 32'h10020874, 32'h00000003, 32'h00000874};
#498 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'had040000, 32'h10020874, 1'b1, 32'h00000003, 32'h00000002, 32'h00000000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10020874, 32'h00000002, 32'h10020874, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020874, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#498 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000000, 32'h00000023, 32'h00f000f0, 32'h10020874, 32'h00000003, 32'h00000002};
#498 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h07c, 10'h000, 12'hfff};
#499 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h00000023, 32'h00f000f0, 32'h10010ffc, 32'h00400024, 32'h00400024};
#499 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h00400024, 32'h00400024, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'h1f, 32'h00400024, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#499 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h07c, 10'h000, 12'hfff};
#500 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00fa00fa, 32'h10010ff8, 32'hxxxxxxxx, 32'h10020874};
#500 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h07d, 10'h000, 12'hfff};
#500 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h10020874, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020874, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#500 bmem_addr <= 'h020d;
#501 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h00000874, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000874, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#501 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00fa00fa, 32'h10010ff4, 32'hxxxxxxxx, 32'h00000874};
#502 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000068, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000068, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#502 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h00fa00fa, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000068};
#503 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#503 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00fa00fa, 32'h10011000, 32'h00000000, 32'h10010ff0};
#504 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400144, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0040, 1'b0, 5'bxxxxx, 1'bx, 32'h00400024, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#504 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00fa00fa, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#504 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h07e, 10'h000, 12'hfff};
#504 bmem_addr <= 'h020e;
#505 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h0c1000d3, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0040, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400028, 32'h000000d3, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#505 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00fa00fa, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#506 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040034c, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10020000, 32'h00000000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#506 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00fa00fa, 32'h10030000, 32'h00000023, 32'h10020000};
#507 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400350, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#507 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00fa00fa, 32'h10030000, 32'h00000023, 32'h00000000};
#508 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h07f, 10'h000, 12'hfff};
#508 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400354, 32'h8c220004, 32'h10030004, 1'b0, 32'h00fa00fa, 32'h00000002, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000002, 32'h10030004, 5'h02, 32'h00fa00fa, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#508 bmem_addr <= 'h020f;
#508 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000023, 32'h00fa00fa, 32'h10030004, 32'h00fa00fa, 32'h00000002};
#509 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400358, 32'h00021402, 32'h000000fa, 1'b0, 32'hxxxxxxxx, 32'h00fa00fa, 32'h00000000, 16'h0040, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00fa00fa, 32'h000000fa, 5'h02, 32'h000000fa, 32'h00001402, 32'h00000010, 32'h00fa00fa, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#509 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00fa00fa, 32'h000000fa, 32'hxxxxxxxx, 32'h00fa00fa};
#510 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040035c, 32'h304201ff, 32'h000000fa, 1'b0, 32'hxxxxxxxx, 32'h000000fa, 32'h00000000, 16'h0040, 1'b1, 5'bx0000, 1'b0, 32'h000000fa, 32'h000000fa, 32'h000000fa, 5'h02, 32'h000000fa, 32'h000001ff, 32'h000000fa, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#510 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00fa00fa, 32'h000000fa, 32'hxxxxxxxx, 32'h000000fa};
#511 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400360, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0040, 1'b0, 5'bxxxxx, 1'bx, 32'h00400028, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#511 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00fa00fa, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#512 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h080, 10'h000, 12'hccc};
#512 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h00022300, 32'h000fa000, 1'b0, 32'h00000023, 32'h000000fa, 32'h00000000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000000fa, 32'h000fa000, 5'h04, 32'h000fa000, 32'h00002300, 32'h0000000c, 32'h000000fa, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#512 smem_addr <= 'h008;
#512 bmem_addr <= 'h0300;
#512 charcode  <= 'h03;
#512 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00fa00fa, 32'h000fa000, 32'h00000023, 32'h000000fa};
#513 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h0c1000de, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0040, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400030, 32'h000000de, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#513 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00fa00fa, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#514 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400378, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10030000, 32'h00000000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#514 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00fa00fa, 32'h10030000, 32'h00000023, 32'h10030000};
#515 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040037c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h00000000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#515 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00fa00fa, 32'h10030000, 32'h00000023, 32'h00000000};
#516 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h081, 10'h000, 12'hccc};
#516 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400380, 32'hac240008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h000fa000, 32'h00000000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h000fa000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#516 bmem_addr <= 'h0301;
#516 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000023, 32'h00fa00fa, 32'h10030008, 32'hxxxxxxxx, 32'h000fa000};
#517 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400384, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000fa000, 16'h0040, 1'b0, 5'bxxxxx, 1'bx, 32'h00400030, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#517 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00fa00fa, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#518 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h0c1000d9, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h000fa000, 16'h0040, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400034, 32'h000000d9, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#518 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h00fa00fa, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#519 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400364, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10030000, 32'h000fa000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#519 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h00fa00fa, 32'h10030000, 32'h00000023, 32'h10030000};
#520 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01040104, 32'h10030000, 32'h00000023, 32'h00000000};
#520 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h082, 10'h000, 12'hccc};
#520 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400368, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h000fa000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#520 bmem_addr <= 'h0302;
#521 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040036c, 32'h8c220004, 32'h10030004, 1'b0, 32'h01040104, 32'h000000fa, 32'h000fa000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h000000fa, 32'h10030004, 5'h02, 32'h01040104, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#521 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000023, 32'h01040104, 32'h10030004, 32'h01040104, 32'h000000fa};
#522 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400370, 32'h304201ff, 32'h00000104, 1'b0, 32'hxxxxxxxx, 32'h01040104, 32'h000fa000, 16'h0040, 1'b1, 5'bx0000, 1'b0, 32'h01040104, 32'h01040104, 32'h00000104, 5'h02, 32'h00000104, 32'h000001ff, 32'h01040104, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#522 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01040104, 32'h00000104, 32'hxxxxxxxx, 32'h01040104};
#523 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400374, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000fa000, 16'h0040, 1'b0, 5'bxxxxx, 1'bx, 32'h00400034, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#523 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h01040104, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#524 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h083, 10'h000, 12'hccc};
#524 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h00021142, 32'h00000008, 1'b0, 32'hxxxxxxxx, 32'h00000104, 32'h000fa000, 16'h0040, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00000104, 32'h00000008, 5'h02, 32'h00000008, 32'h00001142, 32'h00000005, 32'h00000104, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#524 bmem_addr <= 'h0303;
#524 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000023, 32'h01040104, 32'h00000008, 32'hxxxxxxxx, 32'h00000104};
#525 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h24040001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h000fa000, 32'h000fa000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h000fa000, 32'h00000001, 5'h04, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#525 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01040104, 32'h00000001, 32'hxxxxxxxx, 32'h000fa000};
#526 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h00442004, 32'h00000100, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h000fa000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000008, 32'h00000001, 32'h00000100, 5'h04, 32'h00000100, 32'h00002004, 32'h00000008, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#526 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01040104, 32'h00000100, 32'hxxxxxxxx, 32'h00000001};
#527 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h0c1000e6, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h000fa000, 16'h0040, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400044, 32'h000000e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#527 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h01040104, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#528 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400398, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10030000, 32'h000fa000, 16'h0040, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#528 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h084, 10'h000, 12'h999};
#528 bmem_addr <= 'h0304;
#528 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01040104, 32'h10030000, 32'h00000023, 32'h10030000};
#529 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040039c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h000fa000, 16'h0040, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#529 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01040104, 32'h10030000, 32'h00000023, 32'h00000000};
#530 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a0, 32'hac24000c, 32'h1003000c, 1'b1, 32'hxxxxxxxx, 32'h00000100, 32'h000fa000, 16'h0040, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000100, 32'h1003000c, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10030000, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#530 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b1, 32'h00000003, 32'h00000023, 32'h00000023, 32'h01040104, 32'h1003000c, 32'hxxxxxxxx, 32'h00000100};
#531 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a4, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000fa000, 16'h0100, 1'b0, 5'bxxxxx, 1'bx, 32'h00400044, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#531 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h01040104, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#532 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h085, 10'h000, 12'h999};
#532 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h2404000f, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h00000100, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000100, 32'h0000000f, 5'h04, 32'h0000000f, 32'h0000000f, 32'h00000000, 32'h0000000f, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#532 bmem_addr <= 'h0305;
#532 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000023, 32'h01040104, 32'h0000000f, 32'hxxxxxxxx, 32'h00000100};
#533 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h0c100066, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h000fa000, 16'h0100, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h0040004c, 32'h00000066, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#533 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h01040104, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#534 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#534 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h01040104, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#535 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h00400024, 32'h0040004c, 32'h000fa000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#535 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h00000023, 32'h01040104, 32'h10010ffc, 32'h00400024, 32'h0040004c};
#535 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h085, 10'h000, 12'h999};
#536 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h01040104, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#536 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h000fa000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#536 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h086, 10'h000, 12'h999};
#536 bmem_addr <= 'h0306;
#537 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h000fa000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#537 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h01040104, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#538 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h000fa000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#538 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h01040104, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#539 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10030000, 32'h000fa000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#539 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01040104, 32'h10030000, 32'h00000023, 32'h10030000};
#539 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h086, 10'h000, 12'h999};
#540 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h010e010e, 32'h10030000, 32'h00000023, 32'h00000000};
#540 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h087, 10'h000, 12'hf20};
#540 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#540 bmem_addr <= 'h0307;
#541 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8c220000, 32'h10030000, 1'b0, 32'h00000023, 32'h00000008, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000008, 32'h10030000, 5'h02, 32'h00000023, 32'h00000000, 32'h10030000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#541 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h010e010e, 32'h10030000, 32'h00000023, 32'h00000008};
#542 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h1040000f, 32'h00000023, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000fa000, 16'h0100, 1'b0, 5'b1xx01, 1'b0, 32'h00000023, 32'h00000000, 32'h00000023, 5'hxx, 32'hxxxxxxxx, 32'h0000000f, 32'h00000023, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#542 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000043, 32'h00000023, 32'h010e010e, 32'h00000023, 32'hxxxxxxxx, 32'h00000000};
#543 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h00024821, 32'h00000023, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000023, 32'h00000023, 5'h09, 32'h00000023, 32'h00004821, 32'h00000000, 32'h00000023, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#543 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000043, 32'h00000023, 32'h010e010e, 32'h00000023, 32'hxxxxxxxx, 32'h00000023};
#544 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h088, 10'h000, 12'hf20};
#544 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c0, 32'h24020000, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h00000023, 32'h00000000, 5'h02, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#544 bmem_addr <= 'h0308;
#544 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h010e010e, 32'h00000000, 32'hxxxxxxxx, 32'h00000023};
#545 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c4, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10030000, 32'h000fa000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#545 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h010e010e, 32'h10010000, 32'h00000000, 32'h10030000};
#546 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c8, 32'h34280008, 32'h10010008, 1'b0, 32'h0000001c, 32'hxxxxxxxx, 32'h000fa000, 16'h0100, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010008, 5'h08, 32'h10010008, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#546 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000023, 32'h010e010e, 32'h10010008, 32'h0000001c, 32'hxxxxxxxx};
#547 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001cc, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h000fa000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#547 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h010e010e, 32'h10010000, 32'h00000000, 32'h10010000};
#548 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h089, 10'h000, 12'hf20};
#548 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d0, 32'h342a0018, 32'h10010018, 1'b0, 32'h0000003b, 32'hxxxxxxxx, 32'h000fa000, 16'h0100, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010018, 5'h0a, 32'h10010018, 32'h00000018, 32'h10010000, 32'h00000018, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#548 bmem_addr <= 'h0309;
#548 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h00000023, 32'h010e010e, 32'h10010018, 32'h0000003b, 32'hxxxxxxxx};
#549 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d4, 32'h01485022, 32'h00000010, 1'b0, 32'hxxxxxxxx, 32'h10010008, 32'h000fa000, 16'h0100, 1'b1, 5'b1xx01, 1'b0, 32'h10010018, 32'h10010008, 32'h00000010, 5'h0a, 32'h00000010, 32'h00005022, 32'h10010018, 32'h10010008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#549 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h00000023, 32'h010e010e, 32'h00000010, 32'hxxxxxxxx, 32'h10010008};
#550 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h000fa000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#550 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h010e010e, 32'h10010000, 32'h00000000, 32'h10010000};
#551 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#551 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h010e010e, 32'h10010000, 32'h00000000, 32'h00000000};
#552 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h08a, 10'h000, 12'hf20};
#552 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010008, 1'b0, 32'h0000001c, 32'h10010008, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h10010008, 32'h10010008, 5'h08, 32'h0000001c, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#552 bmem_addr <= 'h030a;
#552 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000023, 32'h010e010e, 32'h10010008, 32'h0000001c, 32'h10010008};
#553 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000004, 5'h02, 32'h00000004, 32'h00000004, 32'h00000000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#553 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000023, 32'h010e010e, 32'h00000004, 32'hxxxxxxxx, 32'h00000000};
#554 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'hfffffff9, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000fa000, 16'h0100, 1'b0, 5'b1xx01, 1'b0, 32'h0000001c, 32'h00000023, 32'hfffffff9, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001c, 32'h00000023, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#554 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h010e010e, 32'hfffffff9, 32'hxxxxxxxx, 32'h00000023};
#555 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h000fa000, 16'h0100, 1'b1, 5'b1x011, 1'b0, 32'h00000004, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h00000004, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#555 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h010e010e, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#556 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h08b, 10'h000, 12'hf20};
#556 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000fa000, 16'h0100, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#556 bmem_addr <= 'h030b;
#556 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h010e010e, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#557 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h000fa000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#557 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h010e010e, 32'h10010000, 32'h00000000, 32'h00000001};
#558 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010004, 1'b0, 32'h00000003, 32'h00000004, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000004, 32'h10010004, 5'h01, 32'h10010004, 32'h00000821, 32'h10010000, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#558 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h00000023, 32'h010e010e, 32'h10010004, 32'h00000003, 32'h00000004};
#559 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h1001000c, 1'b0, 32'h00000023, 32'h0000001c, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010004, 32'h0000001c, 32'h1001000c, 5'h08, 32'h00000023, 32'h00000008, 32'h10010004, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#559 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000023, 32'h010e010e, 32'h1001000c, 32'h00000023, 32'h0000001c};
#560 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000023, 32'h01180118, 32'h00000008, 32'hxxxxxxxx, 32'h00000004};
#560 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000008, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000004, 32'h00000004, 32'h00000008, 5'h02, 32'h00000008, 32'h00000004, 32'h00000004, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#560 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h08c, 10'h000, 12'hf20};
#560 bmem_addr <= 'h030c;
#561 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000fa000, 16'h0100, 1'b0, 5'b1xx01, 1'b1, 32'h00000023, 32'h00000023, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h00000023, 32'h00000023, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#561 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01180118, 32'h00000000, 32'hxxxxxxxx, 32'h00000023};
#562 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f8, 32'h00021082, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000008, 32'h000fa000, 16'h0100, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00000008, 32'h00000002, 5'h02, 32'h00000002, 32'h00001082, 32'h00000002, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#562 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01180118, 32'h00000002, 32'hxxxxxxxx, 32'h00000008};
#563 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001fc, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h0040004c, 32'h0040004c, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'h1f, 32'h0040004c, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#563 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h00000023, 32'h01180118, 32'h10010ffc, 32'h0040004c, 32'h0040004c};
#564 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h08d, 10'h000, 12'hf20};
#564 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400200, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000023, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#564 bmem_addr <= 'h030d;
#564 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h01180118, 32'h10010ff8, 32'hxxxxxxxx, 32'h00000023};
#565 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400204, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h00000023, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000023, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#565 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h01180118, 32'h10010ff4, 32'hxxxxxxxx, 32'h00000023};
#566 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400208, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000010, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#566 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h01180118, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000010};
#567 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040020c, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#567 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01180118, 32'h10011000, 32'h00000000, 32'h10010ff0};
#568 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400210, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h000fa000, 16'h0100, 1'b0, 5'bxxxxx, 1'bx, 32'h0040004c, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#568 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h01180118, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#568 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h08e, 10'h000, 12'hf20};
#568 bmem_addr <= 'h030e;
#569 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h00028021, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000002, 5'h10, 32'h00000002, 32'hxxxx8021, 32'h00000000, 32'h00000002, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#569 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01180118, 32'h00000002, 32'hxxxxxxxx, 32'h00000002};
#570 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h0c1000e2, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h000fa000, 16'h0100, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400054, 32'h000000e2, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#570 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h01180118, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#571 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400388, 32'h3c011003, 32'h10030000, 1'b0, 32'h00000023, 32'h10010004, 32'h000fa000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010004, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#571 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01180118, 32'h10030000, 32'h00000023, 32'h10010004};
#572 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040038c, 32'h00200821, 32'h10030000, 1'b0, 32'h00000023, 32'h00000000, 32'h000fa000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#572 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01180118, 32'h10030000, 32'h00000023, 32'h00000000};
#572 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h08f, 10'h000, 12'hf20};
#572 bmem_addr <= 'h030f;
#573 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400390, 32'hac200008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h00000000, 32'h000fa000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#573 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h00000023, 32'h01180118, 32'h10030008, 32'hxxxxxxxx, 32'h00000000};
#574 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400394, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0100, 1'b0, 5'bxxxxx, 1'bx, 32'h00400054, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#574 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h01180118, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#575 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400054, 32'h1200ffef, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0100, 1'b0, 5'b1xx01, 1'b0, 32'h00000002, 32'h00000000, 32'h00000002, 5'hxx, 32'hxxxxxxxx, 32'hffffffef, 32'h00000002, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#575 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01180118, 32'h00000002, 32'hxxxxxxxx, 32'h00000000};
#576 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h090, 10'h000, 12'hf20};
#576 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400058, 32'h20010001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h10030000, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h10030000, 32'h00000001, 5'h01, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#576 smem_addr <= 'h009;
#576 bmem_addr <= 'h0000;
#576 charcode  <= 'h00;
#576 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01180118, 32'h00000001, 32'hxxxxxxxx, 32'h10030000};
#577 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040005c, 32'h14300005, 32'hffffffff, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0100, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000002, 32'hffffffff, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000001, 32'h00000002, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#577 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h00000023, 32'h01180118, 32'hffffffff, 32'hxxxxxxxx, 32'h00000002};
#578 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400074, 32'h20010002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000001, 32'h00000002, 5'h01, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#578 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01180118, 32'h00000002, 32'hxxxxxxxx, 32'h00000001};
#579 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400078, 32'h14300005, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0100, 1'b0, 5'b1xx01, 1'b1, 32'h00000002, 32'h00000002, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000002, 32'h00000002, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#579 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01180118, 32'h00000000, 32'hxxxxxxxx, 32'h00000002};
#580 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h00000023, 32'h01220122, 32'h00000016, 32'hxxxxxxxx, 32'h00000015};
#580 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h091, 10'h000, 12'hf20};
#580 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040007c, 32'h22310001, 32'h00000016, 1'b0, 32'hxxxxxxxx, 32'h00000015, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000015, 32'h00000015, 32'h00000016, 5'h11, 32'h00000016, 32'h00000001, 32'h00000015, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#580 bmem_addr <= 'h0001;
#581 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400080, 32'h2a210028, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0100, 1'b1, 5'b1x011, 1'b0, 32'h00000016, 32'h00000002, 32'h00000001, 5'h01, 32'h00000001, 32'h00000028, 32'h00000016, 32'h00000028, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#581 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01220122, 32'h00000001, 32'hxxxxxxxx, 32'h00000002};
#582 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400084, 32'h1420ffe3, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0100, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hffffffe3, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#582 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01220122, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#583 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h24040002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#583 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01220122, 32'h00000002, 32'hxxxxxxxx, 32'h0000000f};
#584 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00112821, 32'h00000016, 1'b0, 32'hxxxxxxxx, 32'h00000016, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000016, 32'h00000016, 5'h05, 32'h00000016, 32'h00002821, 32'h00000000, 32'h00000016, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#584 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h00000023, 32'h01220122, 32'h00000016, 32'hxxxxxxxx, 32'h00000016};
#584 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h092, 10'h000, 12'hf20};
#584 bmem_addr <= 'h0002;
#585 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h00123021, 32'h0000000d, 1'b0, 32'hxxxxxxxx, 32'h0000000d, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000d, 32'h0000000d, 5'h06, 32'h0000000d, 32'h00003021, 32'h00000000, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#585 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h00000023, 32'h01220122, 32'h0000000d, 32'hxxxxxxxx, 32'h0000000d};
#586 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h0c10003e, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0100, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400024, 32'h0000003e, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#586 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h00000023, 32'h01220122, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#587 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000f8, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#587 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h01220122, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#588 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h0040004c, 32'h00400024, 32'h00000000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#588 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h00000023, 32'h01220122, 32'h10010ffc, 32'h0040004c, 32'h00400024};
#588 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h093, 10'h000, 12'hf20};
#588 bmem_addr <= 'h0003;
#589 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h01220122, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#589 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#590 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#590 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h01220122, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#591 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#591 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000023, 32'h01220122, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#592 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h094, 10'h000, 12'hf20};
#592 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#592 bmem_addr <= 'h0004;
#592 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01220122, 32'h10020000, 32'h00000000, 32'h00000001};
#593 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0100, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'hxxxxxxxx, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#593 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01220122, 32'h10020000, 32'h00000000, 32'hxxxxxxxx};
#594 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h00064940, 32'h000001a0, 1'b0, 32'hxxxxxxxx, 32'h0000000d, 32'h00000000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000d, 32'h000001a0, 5'h09, 32'h000001a0, 32'h00004940, 32'h00000005, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#594 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01220122, 32'h000001a0, 32'hxxxxxxxx, 32'h0000000d};
#595 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h000650c0, 32'h00000068, 1'b0, 32'hxxxxxxxx, 32'h0000000d, 32'h00000000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000d, 32'h00000068, 5'h0a, 32'h00000068, 32'h000050c0, 32'h00000003, 32'h0000000d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#595 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h00000023, 32'h01220122, 32'h00000068, 32'hxxxxxxxx, 32'h0000000d};
#596 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h095, 10'h000, 12'hf20};
#596 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h012a4820, 32'h00000208, 1'b0, 32'hxxxxxxxx, 32'h00000068, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h000001a0, 32'h00000068, 32'h00000208, 5'h09, 32'h00000208, 32'h00004820, 32'h000001a0, 32'h00000068, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#596 bmem_addr <= 'h0005;
#596 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h00000023, 32'h01220122, 32'h00000208, 32'hxxxxxxxx, 32'h00000068};
#597 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h01254820, 32'h0000021e, 1'b0, 32'hxxxxxxxx, 32'h00000016, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000208, 32'h00000016, 32'h0000021e, 5'h09, 32'h0000021e, 32'h00004820, 32'h00000208, 32'h00000016, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#597 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h00000000, 32'h00000023, 32'h01220122, 32'h0000021e, 32'hxxxxxxxx, 32'h00000016};
#598 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h00094880, 32'h00000878, 1'b0, 32'hxxxxxxxx, 32'h0000021e, 32'h00000000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000021e, 32'h00000878, 5'h09, 32'h00000878, 32'h00004880, 32'h00000002, 32'h0000021e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#598 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01220122, 32'h00000878, 32'hxxxxxxxx, 32'h0000021e};
#599 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h01094020, 32'h10020878, 1'b0, 32'h00000000, 32'h00000878, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000878, 32'h10020878, 5'h08, 32'h10020878, 32'h00004020, 32'h10020000, 32'h00000878, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#599 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h00000023, 32'h01220122, 32'h10020878, 32'h00000000, 32'h00000878};
#600 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h012c012c, 32'h10020878, 32'h00000000, 32'h00000002};
#600 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'had040000, 32'h10020878, 1'b1, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10020878, 32'h00000002, 32'h10020878, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020878, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#600 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h096, 10'h000, 12'hf20};
#600 bmem_addr <= 'h0006;
#601 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001b, 32'h012c012c, 32'h10010ffc, 32'h00400024, 32'h00400024};
#601 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h00400024, 32'h00400024, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'h1f, 32'h00400024, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#601 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h096, 10'h000, 12'hf20};
#602 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h10020878, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020878, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#602 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h012c012c, 32'h10010ff8, 32'hxxxxxxxx, 32'h10020878};
#603 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h00000878, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000878, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#603 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h012c012c, 32'h10010ff4, 32'hxxxxxxxx, 32'h00000878};
#604 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000068, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000068, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#604 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h012c012c, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000068};
#604 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h097, 10'h000, 12'hf20};
#604 bmem_addr <= 'h0007;
#605 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#605 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h012c012c, 32'h10011000, 32'h00000000, 32'h10010ff0};
#606 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400144, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0100, 1'b0, 5'bxxxxx, 1'bx, 32'h00400024, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#606 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h012c012c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#607 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h0c1000d3, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0100, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400028, 32'h000000d3, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#607 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h012c012c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#608 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040034c, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001b, 32'h10020000, 32'h00000000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#608 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h098, 10'h000, 12'hf20};
#608 bmem_addr <= 'h0008;
#608 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h012c012c, 32'h10030000, 32'h0000001b, 32'h10020000};
#609 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400350, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000000, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#609 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h012c012c, 32'h10030000, 32'h0000001b, 32'h00000000};
#610 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400354, 32'h8c220004, 32'h10030004, 1'b0, 32'h012c012c, 32'h00000002, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000002, 32'h10030004, 5'h02, 32'h012c012c, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#610 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h012c012c, 32'h10030004, 32'h012c012c, 32'h00000002};
#611 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400358, 32'h00021402, 32'h0000012c, 1'b0, 32'hxxxxxxxx, 32'h012c012c, 32'h00000000, 16'h0100, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h012c012c, 32'h0000012c, 5'h02, 32'h0000012c, 32'h00001402, 32'h00000010, 32'h012c012c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#611 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h012c012c, 32'h0000012c, 32'hxxxxxxxx, 32'h012c012c};
#612 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040035c, 32'h304201ff, 32'h0000012c, 1'b0, 32'hxxxxxxxx, 32'h0000012c, 32'h00000000, 16'h0100, 1'b1, 5'bx0000, 1'b0, 32'h0000012c, 32'h0000012c, 32'h0000012c, 5'h02, 32'h0000012c, 32'h000001ff, 32'h0000012c, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#612 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h012c012c, 32'h0000012c, 32'hxxxxxxxx, 32'h0000012c};
#612 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h099, 10'h000, 12'hf20};
#612 bmem_addr <= 'h0009;
#613 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400360, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0100, 1'b0, 5'bxxxxx, 1'bx, 32'h00400028, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#613 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h012c012c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#614 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h00022300, 32'h0012c000, 1'b0, 32'h00000000, 32'h0000012c, 32'h00000000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000012c, 32'h0012c000, 5'h04, 32'h0012c000, 32'h00002300, 32'h0000000c, 32'h0000012c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#614 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h012c012c, 32'h0012c000, 32'h00000000, 32'h0000012c};
#615 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h0c1000de, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0100, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400030, 32'h000000de, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#615 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h012c012c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#616 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400378, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001b, 32'h10030000, 32'h00000000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#616 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h09a, 10'h000, 12'hf20};
#616 bmem_addr <= 'h000a;
#616 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h012c012c, 32'h10030000, 32'h0000001b, 32'h10030000};
#617 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040037c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000000, 32'h00000000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#617 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h012c012c, 32'h10030000, 32'h0000001b, 32'h00000000};
#618 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400380, 32'hac240008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h0012c000, 32'h00000000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h0012c000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#618 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h012c012c, 32'h10030008, 32'hxxxxxxxx, 32'h0012c000};
#619 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400384, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0012c000, 16'h0100, 1'b0, 5'bxxxxx, 1'bx, 32'h00400030, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#619 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h012c012c, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#620 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01360136, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#620 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h09b, 10'h000, 12'hf20};
#620 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h0c1000d9, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h0012c000, 16'h0100, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400034, 32'h000000d9, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#620 bmem_addr <= 'h000b;
#621 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400364, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001b, 32'h10030000, 32'h0012c000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#621 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01360136, 32'h10030000, 32'h0000001b, 32'h10030000};
#622 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400368, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000000, 32'h0012c000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#622 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01360136, 32'h10030000, 32'h0000001b, 32'h00000000};
#623 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040036c, 32'h8c220004, 32'h10030004, 1'b0, 32'h01360136, 32'h0000012c, 32'h0012c000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h0000012c, 32'h10030004, 5'h02, 32'h01360136, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#623 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h01360136, 32'h10030004, 32'h01360136, 32'h0000012c};
#624 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400370, 32'h304201ff, 32'h00000136, 1'b0, 32'hxxxxxxxx, 32'h01360136, 32'h0012c000, 16'h0100, 1'b1, 5'bx0000, 1'b0, 32'h01360136, 32'h01360136, 32'h00000136, 5'h02, 32'h00000136, 32'h000001ff, 32'h01360136, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#624 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01360136, 32'h00000136, 32'hxxxxxxxx, 32'h01360136};
#624 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h09c, 10'h000, 12'hf20};
#624 bmem_addr <= 'h000c;
#625 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400374, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0012c000, 16'h0100, 1'b0, 5'bxxxxx, 1'bx, 32'h00400034, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#625 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01360136, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#626 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h00021142, 32'h00000009, 1'b0, 32'hxxxxxxxx, 32'h00000136, 32'h0012c000, 16'h0100, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00000136, 32'h00000009, 5'h02, 32'h00000009, 32'h00001142, 32'h00000005, 32'h00000136, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#626 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h01360136, 32'h00000009, 32'hxxxxxxxx, 32'h00000136};
#627 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h24040001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h0012c000, 32'h0012c000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0012c000, 32'h00000001, 5'h04, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#627 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01360136, 32'h00000001, 32'hxxxxxxxx, 32'h0012c000};
#628 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h00442004, 32'h00000200, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h0012c000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000009, 32'h00000001, 32'h00000200, 5'h04, 32'h00000200, 32'h00002004, 32'h00000009, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#628 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000000, 32'h0000001b, 32'h01360136, 32'h00000200, 32'hxxxxxxxx, 32'h00000001};
#628 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h09d, 10'h000, 12'hf20};
#628 bmem_addr <= 'h000d;
#629 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h0c1000e6, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h0012c000, 16'h0100, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h00400044, 32'h000000e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#629 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01360136, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#630 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400398, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001b, 32'h10030000, 32'h0012c000, 16'h0100, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#630 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01360136, 32'h10030000, 32'h0000001b, 32'h10030000};
#631 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040039c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000000, 32'h0012c000, 16'h0100, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#631 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01360136, 32'h10030000, 32'h0000001b, 32'h00000000};
#632 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h09e, 10'h000, 12'hf20};
#632 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a0, 32'hac24000c, 32'h1003000c, 1'b1, 32'hxxxxxxxx, 32'h00000200, 32'h0012c000, 16'h0100, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000200, 32'h1003000c, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10030000, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#632 bmem_addr <= 'h000e;
#632 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b1, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h01360136, 32'h1003000c, 32'hxxxxxxxx, 32'h00000200};
#633 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a4, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0012c000, 16'h0200, 1'b0, 5'bxxxxx, 1'bx, 32'h00400044, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#633 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01360136, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#634 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h2404000f, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h00000200, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000200, 32'h0000000f, 5'h04, 32'h0000000f, 32'h0000000f, 32'h00000000, 32'h0000000f, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#634 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h01360136, 32'h0000000f, 32'hxxxxxxxx, 32'h00000200};
#635 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h0c100066, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h0012c000, 16'h0200, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000002, 32'hxxxxxxxx, 5'h1f, 32'h0040004c, 32'h00000066, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#635 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01360136, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000002};
#636 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#636 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h09f, 10'h000, 12'hf20};
#636 bmem_addr <= 'h000f;
#636 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01360136, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#637 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h00400024, 32'h0040004c, 32'h0012c000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#637 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001b, 32'h01360136, 32'h10010ffc, 32'h00400024, 32'h0040004c};
#637 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h09f, 10'h000, 12'hf20};
#638 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01360136, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#638 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0012c000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#639 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0012c000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#639 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01360136, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#640 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01400140, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#640 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0a0, 10'h000, 12'hf20};
#640 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h0012c000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#640 smem_addr <= 'h00a;
#640 bmem_addr <= 'h0000;
#641 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001b, 32'h10030000, 32'h0012c000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#641 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h10030000, 32'h0000001b, 32'h10030000};
#641 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0a0, 10'h000, 12'hf20};
#642 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000000, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#642 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h10030000, 32'h0000001b, 32'h00000000};
#643 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8c220000, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000009, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000009, 32'h10030000, 5'h02, 32'h0000001b, 32'h00000000, 32'h10030000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#643 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h10030000, 32'h0000001b, 32'h00000009};
#644 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h1040000f, 32'h0000001b, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0012c000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h0000001b, 32'h00000000, 32'h0000001b, 5'hxx, 32'hxxxxxxxx, 32'h0000000f, 32'h0000001b, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#644 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h0000001b, 32'h01400140, 32'h0000001b, 32'hxxxxxxxx, 32'h00000000};
#644 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0a1, 10'h000, 12'hf20};
#644 bmem_addr <= 'h0001;
#645 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h00024821, 32'h0000001b, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000001b, 32'h0000001b, 5'h09, 32'h0000001b, 32'h00004821, 32'h00000000, 32'h0000001b, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#645 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h0000001b, 32'h01400140, 32'h0000001b, 32'hxxxxxxxx, 32'h0000001b};
#646 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c0, 32'h24020000, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h0000001b, 32'h00000000, 5'h02, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#646 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b};
#647 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c4, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10030000, 32'h0012c000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#647 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h10010000, 32'h00000000, 32'h10030000};
#648 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c8, 32'h34280008, 32'h10010008, 1'b0, 32'h0000001c, 32'hxxxxxxxx, 32'h0012c000, 16'h0200, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010008, 5'h08, 32'h10010008, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#648 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h01400140, 32'h10010008, 32'h0000001c, 32'hxxxxxxxx};
#648 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0a2, 10'h000, 12'hf20};
#648 bmem_addr <= 'h0002;
#649 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001cc, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h0012c000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#649 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h10010000, 32'h00000000, 32'h10010000};
#650 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d0, 32'h342a0018, 32'h10010018, 1'b0, 32'h0000003b, 32'hxxxxxxxx, 32'h0012c000, 16'h0200, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010018, 5'h0a, 32'h10010018, 32'h00000018, 32'h10010000, 32'h00000018, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#650 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h0000001b, 32'h01400140, 32'h10010018, 32'h0000003b, 32'hxxxxxxxx};
#651 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d4, 32'h01485022, 32'h00000010, 1'b0, 32'hxxxxxxxx, 32'h10010008, 32'h0012c000, 16'h0200, 1'b1, 5'b1xx01, 1'b0, 32'h10010018, 32'h10010008, 32'h00000010, 5'h0a, 32'h00000010, 32'h00005022, 32'h10010018, 32'h10010008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#651 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001b, 32'h01400140, 32'h00000010, 32'hxxxxxxxx, 32'h10010008};
#652 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h0012c000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#652 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h10010000, 32'h00000000, 32'h10010000};
#652 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0a3, 10'h000, 12'hf20};
#652 bmem_addr <= 'h0003;
#653 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#653 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h10010000, 32'h00000000, 32'h00000000};
#654 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010008, 1'b0, 32'h0000001c, 32'h10010008, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h10010008, 32'h10010008, 5'h08, 32'h0000001c, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#654 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h01400140, 32'h10010008, 32'h0000001c, 32'h10010008};
#655 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000004, 5'h02, 32'h00000004, 32'h00000004, 32'h00000000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#655 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h01400140, 32'h00000004, 32'hxxxxxxxx, 32'h00000000};
#656 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h0012c000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h0000001c, 32'h0000001b, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001c, 32'h0000001b, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#656 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h00000001, 32'hxxxxxxxx, 32'h0000001b};
#656 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0a4, 10'h000, 12'hf20};
#656 bmem_addr <= 'h0004;
#657 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0012c000, 16'h0200, 1'b1, 5'b1x011, 1'b0, 32'h00000004, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h00000004, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#657 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#658 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0012c000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#658 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#659 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h0012c000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#659 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01400140, 32'h10010000, 32'h00000000, 32'h00000001};
#660 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h014a014a, 32'h10010004, 32'h00000003, 32'h00000004};
#660 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010004, 1'b0, 32'h00000003, 32'h00000004, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000004, 32'h10010004, 5'h01, 32'h10010004, 32'h00000821, 32'h10010000, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#660 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0a5, 10'h000, 12'hf20};
#660 bmem_addr <= 'h0005;
#661 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h1001000c, 1'b0, 32'h00000023, 32'h0000001c, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010004, 32'h0000001c, 32'h1001000c, 5'h08, 32'h00000023, 32'h00000008, 32'h10010004, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#661 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h014a014a, 32'h1001000c, 32'h00000023, 32'h0000001c};
#662 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000008, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000004, 32'h00000004, 32'h00000008, 5'h02, 32'h00000008, 32'h00000004, 32'h00000004, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#662 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h014a014a, 32'h00000008, 32'hxxxxxxxx, 32'h00000004};
#663 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000008, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h0012c000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h00000023, 32'h0000001b, 32'h00000008, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h00000023, 32'h0000001b, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#663 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h014a014a, 32'h00000008, 32'hxxxxxxxx, 32'h0000001b};
#664 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0a6, 10'h000, 12'hf20};
#664 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0012c000, 16'h0200, 1'b1, 5'b1x011, 1'b0, 32'h00000008, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h00000008, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#664 bmem_addr <= 'h0006;
#664 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h014a014a, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#665 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0012c000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#665 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h014a014a, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#666 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h0012c000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#666 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h014a014a, 32'h10010000, 32'h00000000, 32'h00000001};
#667 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010008, 1'b0, 32'h0000001c, 32'h00000008, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000008, 32'h10010008, 5'h01, 32'h10010008, 32'h00000821, 32'h10010000, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#667 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h014a014a, 32'h10010008, 32'h0000001c, 32'h00000008};
#668 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010010, 1'b0, 32'h0000001d, 32'h00000023, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010008, 32'h00000023, 32'h10010010, 5'h08, 32'h0000001d, 32'h00000008, 32'h10010008, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#668 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001b, 32'h014a014a, 32'h10010010, 32'h0000001d, 32'h00000023};
#668 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0a7, 10'h000, 12'hf20};
#668 bmem_addr <= 'h0007;
#669 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h0000000c, 1'b0, 32'hxxxxxxxx, 32'h00000008, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000008, 32'h00000008, 32'h0000000c, 5'h02, 32'h0000000c, 32'h00000004, 32'h00000008, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#669 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h014a014a, 32'h0000000c, 32'hxxxxxxxx, 32'h00000008};
#670 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h0012c000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h0000001d, 32'h0000001b, 32'h00000002, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001d, 32'h0000001b, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#670 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h014a014a, 32'h00000002, 32'hxxxxxxxx, 32'h0000001b};
#671 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0012c000, 16'h0200, 1'b1, 5'b1x011, 1'b0, 32'h0000000c, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h0000000c, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#671 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h014a014a, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#672 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0a8, 10'h000, 12'hf20};
#672 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0012c000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#672 bmem_addr <= 'h0008;
#672 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h014a014a, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#673 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h0012c000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#673 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h014a014a, 32'h10010000, 32'h00000000, 32'h00000001};
#674 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h1001000c, 1'b0, 32'h00000023, 32'h0000000c, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h0000000c, 32'h1001000c, 5'h01, 32'h1001000c, 32'h00000821, 32'h10010000, 32'h0000000c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#674 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h014a014a, 32'h1001000c, 32'h00000023, 32'h0000000c};
#675 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010014, 1'b0, 32'h0000001b, 32'h0000001d, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h1001000c, 32'h0000001d, 32'h10010014, 5'h08, 32'h0000001b, 32'h00000008, 32'h1001000c, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#675 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h0000001b, 32'h014a014a, 32'h10010014, 32'h0000001b, 32'h0000001d};
#676 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000010, 1'b0, 32'hxxxxxxxx, 32'h0000000c, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h0000000c, 32'h0000000c, 32'h00000010, 5'h02, 32'h00000010, 32'h00000004, 32'h0000000c, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#676 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001b, 32'h014a014a, 32'h00000010, 32'hxxxxxxxx, 32'h0000000c};
#676 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0a9, 10'h000, 12'hf20};
#676 bmem_addr <= 'h0009;
#677 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h0012c000, 16'h0200, 1'b0, 5'b1xx01, 1'b1, 32'h0000001b, 32'h0000001b, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001b, 32'h0000001b, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#677 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h014a014a, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b};
#678 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f8, 32'h00021082, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0012c000, 16'h0200, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00000010, 32'h00000004, 5'h02, 32'h00000004, 32'h00001082, 32'h00000002, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#678 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h014a014a, 32'h00000004, 32'hxxxxxxxx, 32'h00000010};
#679 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001fc, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h0040004c, 32'h0040004c, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'h1f, 32'h0040004c, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#679 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h0000001b, 32'h014a014a, 32'h10010ffc, 32'h0040004c, 32'h0040004c};
#680 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01540154, 32'h10010ff8, 32'hxxxxxxxx, 32'h0000001b};
#680 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0aa, 10'h000, 12'hf20};
#680 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400200, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001b, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#680 bmem_addr <= 'h000a;
#681 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400204, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001b, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#681 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01540154, 32'h10010ff4, 32'hxxxxxxxx, 32'h0000001b};
#682 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400208, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000010, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#682 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01540154, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000010};
#683 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040020c, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#683 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01540154, 32'h10011000, 32'h00000000, 32'h10010ff0};
#684 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400210, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h0012c000, 16'h0200, 1'b0, 5'bxxxxx, 1'bx, 32'h0040004c, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#684 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01540154, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#684 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0ab, 10'h000, 12'hf20};
#684 bmem_addr <= 'h000b;
#685 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h00028021, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000004, 32'h00000004, 5'h10, 32'h00000004, 32'hxxxx8021, 32'h00000000, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#685 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h01540154, 32'h00000004, 32'hxxxxxxxx, 32'h00000004};
#686 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h0c1000e2, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h0012c000, 16'h0200, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400054, 32'h000000e2, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#686 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01540154, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#687 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400388, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001b, 32'h1001000c, 32'h0012c000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h1001000c, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#687 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01540154, 32'h10030000, 32'h0000001b, 32'h1001000c};
#688 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040038c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000000, 32'h0012c000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#688 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01540154, 32'h10030000, 32'h0000001b, 32'h00000000};
#688 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0ac, 10'h000, 12'hf20};
#688 bmem_addr <= 'h000c;
#689 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400390, 32'hac200008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h00000000, 32'h0012c000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#689 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h01540154, 32'h10030008, 32'hxxxxxxxx, 32'h00000000};
#690 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400394, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0200, 1'b0, 5'bxxxxx, 1'bx, 32'h00400054, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#690 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01540154, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#691 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400054, 32'h1200ffef, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h00000004, 32'h00000000, 32'h00000004, 5'hxx, 32'hxxxxxxxx, 32'hffffffef, 32'h00000004, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#691 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h01540154, 32'h00000004, 32'hxxxxxxxx, 32'h00000000};
#692 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0ad, 10'h000, 12'hf20};
#692 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400058, 32'h20010001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h10030000, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h10030000, 32'h00000001, 5'h01, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#692 bmem_addr <= 'h000d;
#692 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01540154, 32'h00000001, 32'hxxxxxxxx, 32'h10030000};
#693 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040005c, 32'h14300005, 32'hfffffffd, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000004, 32'hfffffffd, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000001, 32'h00000004, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#693 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001b, 32'h01540154, 32'hfffffffd, 32'hxxxxxxxx, 32'h00000004};
#694 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400074, 32'h20010002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000001, 32'h00000002, 5'h01, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#694 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01540154, 32'h00000002, 32'hxxxxxxxx, 32'h00000001};
#695 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400078, 32'h14300005, 32'hfffffffe, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h00000002, 32'h00000004, 32'hfffffffe, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000002, 32'h00000004, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#695 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001b, 32'h01540154, 32'hfffffffe, 32'hxxxxxxxx, 32'h00000004};
#696 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0ae, 10'h000, 12'hf20};
#696 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400090, 32'h20010003, 32'h00000003, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000003, 5'h01, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#696 bmem_addr <= 'h000e;
#696 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01540154, 32'h00000003, 32'hxxxxxxxx, 32'h00000002};
#697 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400094, 32'h14300005, 32'hffffffff, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h00000003, 32'h00000004, 32'hffffffff, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000003, 32'h00000004, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#697 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001b, 32'h01540154, 32'hffffffff, 32'hxxxxxxxx, 32'h00000004};
#698 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ac, 32'h20010004, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000004, 5'h01, 32'h00000004, 32'h00000004, 32'h00000000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#698 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h01540154, 32'h00000004, 32'hxxxxxxxx, 32'h00000003};
#699 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000b0, 32'h1430ffd8, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0200, 1'b0, 5'b1xx01, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'hffffffd8, 32'h00000004, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#699 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01540154, 32'h00000000, 32'hxxxxxxxx, 32'h00000004};
#700 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h015e015e, 32'h0000000e, 32'hxxxxxxxx, 32'h0000000d};
#700 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0af, 10'h000, 12'hf20};
#700 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000b4, 32'h22520001, 32'h0000000e, 1'b0, 32'hxxxxxxxx, 32'h0000000d, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h0000000d, 32'h0000000d, 32'h0000000e, 5'h12, 32'h0000000e, 32'h00000001, 32'h0000000d, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#700 bmem_addr <= 'h000f;
#701 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000b8, 32'h2a41001e, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0200, 1'b1, 5'b1x011, 1'b0, 32'h0000000e, 32'h00000004, 32'h00000001, 5'h01, 32'h00000001, 32'h0000001e, 32'h0000000e, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#701 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h015e015e, 32'h00000001, 32'hxxxxxxxx, 32'h00000004};
#702 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000bc, 32'h1420ffd5, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0200, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hffffffd5, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#702 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h015e015e, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#703 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h24040002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#703 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h015e015e, 32'h00000002, 32'hxxxxxxxx, 32'h0000000f};
#704 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00112821, 32'h00000016, 1'b0, 32'hxxxxxxxx, 32'h00000016, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000016, 32'h00000016, 5'h05, 32'h00000016, 32'h00002821, 32'h00000000, 32'h00000016, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#704 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h0000001b, 32'h015e015e, 32'h00000016, 32'hxxxxxxxx, 32'h00000016};
#704 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0b0, 10'h000, 12'h0f0};
#704 smem_addr <= 'h00b;
#704 bmem_addr <= 'h0100;
#704 charcode  <= 'h01;
#705 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h00123021, 32'h0000000e, 1'b0, 32'hxxxxxxxx, 32'h0000000e, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000e, 32'h0000000e, 5'h06, 32'h0000000e, 32'h00003021, 32'h00000000, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#705 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h015e015e, 32'h0000000e, 32'hxxxxxxxx, 32'h0000000e};
#706 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h0c10003e, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0200, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400024, 32'h0000003e, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#706 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h015e015e, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#707 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000f8, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#707 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h015e015e, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#708 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h0040004c, 32'h00400024, 32'h00000000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#708 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h0000001b, 32'h015e015e, 32'h10010ffc, 32'h0040004c, 32'h00400024};
#708 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0b1, 10'h000, 12'h0f0};
#708 bmem_addr <= 'h0101;
#709 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h015e015e, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#709 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#710 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#710 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h015e015e, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#711 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#711 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h015e015e, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#712 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0b2, 10'h000, 12'h0f0};
#712 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#712 bmem_addr <= 'h0102;
#712 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h015e015e, 32'h10020000, 32'h00000000, 32'h00000001};
#713 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0200, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'hxxxxxxxx, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#713 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h015e015e, 32'h10020000, 32'h00000000, 32'hxxxxxxxx};
#714 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h00064940, 32'h000001c0, 1'b0, 32'hxxxxxxxx, 32'h0000000e, 32'h00000000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000e, 32'h000001c0, 5'h09, 32'h000001c0, 32'h00004940, 32'h00000005, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#714 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h015e015e, 32'h000001c0, 32'hxxxxxxxx, 32'h0000000e};
#715 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h000650c0, 32'h00000070, 1'b0, 32'hxxxxxxxx, 32'h0000000e, 32'h00000000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000e, 32'h00000070, 5'h0a, 32'h00000070, 32'h000050c0, 32'h00000003, 32'h0000000e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#715 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000000, 32'h0000001b, 32'h015e015e, 32'h00000070, 32'hxxxxxxxx, 32'h0000000e};
#716 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0b3, 10'h000, 12'h0f0};
#716 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h012a4820, 32'h00000230, 1'b0, 32'hxxxxxxxx, 32'h00000070, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h000001c0, 32'h00000070, 32'h00000230, 5'h09, 32'h00000230, 32'h00004820, 32'h000001c0, 32'h00000070, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#716 bmem_addr <= 'h0103;
#716 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h015e015e, 32'h00000230, 32'hxxxxxxxx, 32'h00000070};
#717 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h01254820, 32'h00000246, 1'b0, 32'hxxxxxxxx, 32'h00000016, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000230, 32'h00000016, 32'h00000246, 5'h09, 32'h00000246, 32'h00004820, 32'h00000230, 32'h00000016, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#717 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h015e015e, 32'h00000246, 32'hxxxxxxxx, 32'h00000016};
#718 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h00094880, 32'h00000918, 1'b0, 32'hxxxxxxxx, 32'h00000246, 32'h00000000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000246, 32'h00000918, 5'h09, 32'h00000918, 32'h00004880, 32'h00000002, 32'h00000246, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#718 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h015e015e, 32'h00000918, 32'hxxxxxxxx, 32'h00000246};
#719 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h01094020, 32'h10020918, 1'b0, 32'h00000000, 32'h00000918, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h00000918, 32'h10020918, 5'h08, 32'h10020918, 32'h00004020, 32'h10020000, 32'h00000918, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#719 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h015e015e, 32'h10020918, 32'h00000000, 32'h00000918};
#720 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01680168, 32'h10020918, 32'h00000000, 32'h00000002};
#720 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'had040000, 32'h10020918, 1'b1, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10020918, 32'h00000002, 32'h10020918, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10020918, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#720 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b1, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0b4, 10'h000, 12'h0f0};
#720 bmem_addr <= 'h0104;
#721 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001b, 32'h01680168, 32'h10010ffc, 32'h00400024, 32'h00400024};
#721 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h00400024, 32'h00400024, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'h1f, 32'h00400024, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#721 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0b4, 10'h000, 12'h0f0};
#722 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h10020918, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10020918, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#722 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01680168, 32'h10010ff8, 32'hxxxxxxxx, 32'h10020918};
#723 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h00000918, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000918, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#723 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01680168, 32'h10010ff4, 32'hxxxxxxxx, 32'h00000918};
#724 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000070, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000070, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#724 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01680168, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000070};
#724 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0b5, 10'h000, 12'h0f0};
#724 bmem_addr <= 'h0105;
#725 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#725 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01680168, 32'h10011000, 32'h00000000, 32'h10010ff0};
#726 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400144, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0200, 1'b0, 5'bxxxxx, 1'bx, 32'h00400024, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#726 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01680168, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#727 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h0c1000d3, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0200, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400028, 32'h000000d3, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#727 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01680168, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#728 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040034c, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001b, 32'h10020000, 32'h00000000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#728 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0b6, 10'h000, 12'h0f0};
#728 bmem_addr <= 'h0106;
#728 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01680168, 32'h10030000, 32'h0000001b, 32'h10020000};
#729 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400350, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000000, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#729 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01680168, 32'h10030000, 32'h0000001b, 32'h00000000};
#730 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400354, 32'h8c220004, 32'h10030004, 1'b0, 32'h01680168, 32'h00000004, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000004, 32'h10030004, 5'h02, 32'h01680168, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#730 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h01680168, 32'h10030004, 32'h01680168, 32'h00000004};
#731 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400358, 32'h00021402, 32'h00000168, 1'b0, 32'hxxxxxxxx, 32'h01680168, 32'h00000000, 16'h0200, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h01680168, 32'h00000168, 5'h02, 32'h00000168, 32'h00001402, 32'h00000010, 32'h01680168, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#731 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01680168, 32'h00000168, 32'hxxxxxxxx, 32'h01680168};
#732 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040035c, 32'h304201ff, 32'h00000168, 1'b0, 32'hxxxxxxxx, 32'h00000168, 32'h00000000, 16'h0200, 1'b1, 5'bx0000, 1'b0, 32'h00000168, 32'h00000168, 32'h00000168, 5'h02, 32'h00000168, 32'h000001ff, 32'h00000168, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#732 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01680168, 32'h00000168, 32'hxxxxxxxx, 32'h00000168};
#732 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0b7, 10'h000, 12'h0f0};
#732 bmem_addr <= 'h0107;
#733 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400360, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0200, 1'b0, 5'bxxxxx, 1'bx, 32'h00400028, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#733 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01680168, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#734 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h00022300, 32'h00168000, 1'b0, 32'h00000000, 32'h00000168, 32'h00000000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000168, 32'h00168000, 5'h04, 32'h00168000, 32'h00002300, 32'h0000000c, 32'h00000168, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#734 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01680168, 32'h00168000, 32'h00000000, 32'h00000168};
#735 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h0c1000de, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0200, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400030, 32'h000000de, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#735 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01680168, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#736 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400378, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001b, 32'h10030000, 32'h00000000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#736 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0b8, 10'h000, 12'h0f0};
#736 bmem_addr <= 'h0108;
#736 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01680168, 32'h10030000, 32'h0000001b, 32'h10030000};
#737 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040037c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000000, 32'h00000000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#737 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01680168, 32'h10030000, 32'h0000001b, 32'h00000000};
#738 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400380, 32'hac240008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h00168000, 32'h00000000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00168000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#738 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h01680168, 32'h10030008, 32'hxxxxxxxx, 32'h00168000};
#739 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400384, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00168000, 16'h0200, 1'b0, 5'bxxxxx, 1'bx, 32'h00400030, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#739 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01680168, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#740 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01720172, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#740 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0b9, 10'h000, 12'h0f0};
#740 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h0c1000d9, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00168000, 16'h0200, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400034, 32'h000000d9, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#740 bmem_addr <= 'h0109;
#741 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400364, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001b, 32'h10030000, 32'h00168000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#741 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01720172, 32'h10030000, 32'h0000001b, 32'h10030000};
#742 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400368, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000000, 32'h00168000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#742 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01720172, 32'h10030000, 32'h0000001b, 32'h00000000};
#743 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040036c, 32'h8c220004, 32'h10030004, 1'b0, 32'h01720172, 32'h00000168, 32'h00168000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000168, 32'h10030004, 5'h02, 32'h01720172, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#743 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h01720172, 32'h10030004, 32'h01720172, 32'h00000168};
#744 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400370, 32'h304201ff, 32'h00000172, 1'b0, 32'hxxxxxxxx, 32'h01720172, 32'h00168000, 16'h0200, 1'b1, 5'bx0000, 1'b0, 32'h01720172, 32'h01720172, 32'h00000172, 5'h02, 32'h00000172, 32'h000001ff, 32'h01720172, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#744 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01720172, 32'h00000172, 32'hxxxxxxxx, 32'h01720172};
#744 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0ba, 10'h000, 12'h0f0};
#744 bmem_addr <= 'h010a;
#745 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400374, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00168000, 16'h0200, 1'b0, 5'bxxxxx, 1'bx, 32'h00400034, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#745 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01720172, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#746 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h00021142, 32'h0000000b, 1'b0, 32'hxxxxxxxx, 32'h00000172, 32'h00168000, 16'h0200, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00000172, 32'h0000000b, 5'h02, 32'h0000000b, 32'h00001142, 32'h00000005, 32'h00000172, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#746 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h01720172, 32'h0000000b, 32'hxxxxxxxx, 32'h00000172};
#747 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h24040001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00168000, 32'h00168000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00168000, 32'h00000001, 5'h04, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#747 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01720172, 32'h00000001, 32'hxxxxxxxx, 32'h00168000};
#748 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h00442004, 32'h00000800, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00168000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h0000000b, 32'h00000001, 32'h00000800, 5'h04, 32'h00000800, 32'h00002004, 32'h0000000b, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#748 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01720172, 32'h00000800, 32'hxxxxxxxx, 32'h00000001};
#748 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0bb, 10'h000, 12'h0f0};
#748 bmem_addr <= 'h010b;
#749 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h0c1000e6, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00168000, 16'h0200, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400044, 32'h000000e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#749 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01720172, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#750 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400398, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001b, 32'h10030000, 32'h00168000, 16'h0200, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#750 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01720172, 32'h10030000, 32'h0000001b, 32'h10030000};
#751 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040039c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000000, 32'h00168000, 16'h0200, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#751 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01720172, 32'h10030000, 32'h0000001b, 32'h00000000};
#752 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0bc, 10'h000, 12'h0f0};
#752 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a0, 32'hac24000c, 32'h1003000c, 1'b1, 32'hxxxxxxxx, 32'h00000800, 32'h00168000, 16'h0200, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000800, 32'h1003000c, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10030000, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#752 bmem_addr <= 'h010c;
#752 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b1, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h01720172, 32'h1003000c, 32'hxxxxxxxx, 32'h00000800};
#753 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a4, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00168000, 16'h0800, 1'b0, 5'bxxxxx, 1'bx, 32'h00400044, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#753 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01720172, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#754 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h2404000f, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h00000800, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000800, 32'h0000000f, 5'h04, 32'h0000000f, 32'h0000000f, 32'h00000000, 32'h0000000f, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#754 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h01720172, 32'h0000000f, 32'hxxxxxxxx, 32'h00000800};
#755 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h0c100066, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00168000, 16'h0800, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h0040004c, 32'h00000066, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#755 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001b, 32'h01720172, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#756 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#756 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0bd, 10'h000, 12'h0f0};
#756 bmem_addr <= 'h010d;
#756 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01720172, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#757 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h00400024, 32'h0040004c, 32'h00168000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#757 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001b, 32'h01720172, 32'h10010ffc, 32'h00400024, 32'h0040004c};
#757 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0bd, 10'h000, 12'h0f0};
#758 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01720172, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#758 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00168000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#759 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00168000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#759 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h01720172, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#760 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b, 32'h017c017c, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#760 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0be, 10'h000, 12'h0f0};
#760 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00168000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#760 bmem_addr <= 'h010e;
#761 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001b, 32'h10030000, 32'h00168000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#761 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h10030000, 32'h0000001b, 32'h10030000};
#761 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0be, 10'h000, 12'h0f0};
#762 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001b, 32'h00000000, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#762 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h10030000, 32'h0000001b, 32'h00000000};
#763 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8c220000, 32'h10030000, 1'b0, 32'h0000001b, 32'h0000000b, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h0000000b, 32'h10030000, 5'h02, 32'h0000001b, 32'h00000000, 32'h10030000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#763 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h10030000, 32'h0000001b, 32'h0000000b};
#764 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h1040000f, 32'h0000001b, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00168000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h0000001b, 32'h00000000, 32'h0000001b, 5'hxx, 32'hxxxxxxxx, 32'h0000000f, 32'h0000001b, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#764 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h0000001b, 32'h017c017c, 32'h0000001b, 32'hxxxxxxxx, 32'h00000000};
#764 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h0, 4'hf, 4'h0, 10'h0bf, 10'h000, 12'h0f0};
#764 bmem_addr <= 'h010f;
#765 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h00024821, 32'h0000001b, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000001b, 32'h0000001b, 5'h09, 32'h0000001b, 32'h00004821, 32'h00000000, 32'h0000001b, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#765 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h0000001b, 32'h017c017c, 32'h0000001b, 32'hxxxxxxxx, 32'h0000001b};
#766 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c0, 32'h24020000, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h0000001b, 32'h00000000, 5'h02, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#766 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b};
#767 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c4, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10030000, 32'h00168000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#767 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h10010000, 32'h00000000, 32'h10030000};
#768 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c8, 32'h34280008, 32'h10010008, 1'b0, 32'h0000001c, 32'hxxxxxxxx, 32'h00168000, 16'h0800, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010008, 5'h08, 32'h10010008, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#768 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h017c017c, 32'h10010008, 32'h0000001c, 32'hxxxxxxxx};
#768 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0c0, 10'h000, 12'hfff};
#768 smem_addr <= 'h00c;
#768 bmem_addr <= 'h0200;
#768 charcode  <= 'h02;
#769 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001cc, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h00168000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#769 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h10010000, 32'h00000000, 32'h10010000};
#770 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d0, 32'h342a0018, 32'h10010018, 1'b0, 32'h0000003b, 32'hxxxxxxxx, 32'h00168000, 16'h0800, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010018, 5'h0a, 32'h10010018, 32'h00000018, 32'h10010000, 32'h00000018, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#770 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h0000001b, 32'h017c017c, 32'h10010018, 32'h0000003b, 32'hxxxxxxxx};
#771 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d4, 32'h01485022, 32'h00000010, 1'b0, 32'hxxxxxxxx, 32'h10010008, 32'h00168000, 16'h0800, 1'b1, 5'b1xx01, 1'b0, 32'h10010018, 32'h10010008, 32'h00000010, 5'h0a, 32'h00000010, 32'h00005022, 32'h10010018, 32'h10010008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#771 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001b, 32'h017c017c, 32'h00000010, 32'hxxxxxxxx, 32'h10010008};
#772 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h00168000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#772 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h10010000, 32'h00000000, 32'h10010000};
#772 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0c1, 10'h000, 12'hfff};
#772 bmem_addr <= 'h0201;
#773 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#773 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h10010000, 32'h00000000, 32'h00000000};
#774 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010008, 1'b0, 32'h0000001c, 32'h10010008, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h10010008, 32'h10010008, 5'h08, 32'h0000001c, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#774 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h017c017c, 32'h10010008, 32'h0000001c, 32'h10010008};
#775 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000004, 5'h02, 32'h00000004, 32'h00000004, 32'h00000000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#775 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h017c017c, 32'h00000004, 32'hxxxxxxxx, 32'h00000000};
#776 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h00168000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h0000001c, 32'h0000001b, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001c, 32'h0000001b, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#776 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h00000001, 32'hxxxxxxxx, 32'h0000001b};
#776 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0c2, 10'h000, 12'hfff};
#776 bmem_addr <= 'h0202;
#777 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h00168000, 16'h0800, 1'b1, 5'b1x011, 1'b0, 32'h00000004, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h00000004, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#777 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#778 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00168000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#778 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#779 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h00168000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#779 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h017c017c, 32'h10010000, 32'h00000000, 32'h00000001};
#780 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h01860186, 32'h10010004, 32'h00000003, 32'h00000004};
#780 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010004, 1'b0, 32'h00000003, 32'h00000004, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000004, 32'h10010004, 5'h01, 32'h10010004, 32'h00000821, 32'h10010000, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#780 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0c3, 10'h000, 12'hfff};
#780 bmem_addr <= 'h0203;
#781 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h1001000c, 1'b0, 32'h00000023, 32'h0000001c, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010004, 32'h0000001c, 32'h1001000c, 5'h08, 32'h00000023, 32'h00000008, 32'h10010004, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#781 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h01860186, 32'h1001000c, 32'h00000023, 32'h0000001c};
#782 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000008, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000004, 32'h00000004, 32'h00000008, 5'h02, 32'h00000008, 32'h00000004, 32'h00000004, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#782 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h01860186, 32'h00000008, 32'hxxxxxxxx, 32'h00000004};
#783 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000008, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h00168000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h00000023, 32'h0000001b, 32'h00000008, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h00000023, 32'h0000001b, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#783 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h01860186, 32'h00000008, 32'hxxxxxxxx, 32'h0000001b};
#784 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hd, 4'hc, 10'h0c4, 10'h000, 12'hfdc};
#784 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h00168000, 16'h0800, 1'b1, 5'b1x011, 1'b0, 32'h00000008, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h00000008, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#784 bmem_addr <= 'h0204;
#784 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01860186, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#785 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00168000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#785 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01860186, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#786 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h00168000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#786 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01860186, 32'h10010000, 32'h00000000, 32'h00000001};
#787 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010008, 1'b0, 32'h0000001c, 32'h00000008, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000008, 32'h10010008, 5'h01, 32'h10010008, 32'h00000821, 32'h10010000, 32'h00000008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#787 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001b, 32'h01860186, 32'h10010008, 32'h0000001c, 32'h00000008};
#788 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010010, 1'b0, 32'h0000001d, 32'h00000023, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010008, 32'h00000023, 32'h10010010, 5'h08, 32'h0000001d, 32'h00000008, 32'h10010008, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#788 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001b, 32'h01860186, 32'h10010010, 32'h0000001d, 32'h00000023};
#788 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h8, 10'h0c5, 10'h000, 12'hfc8};
#788 bmem_addr <= 'h0205;
#789 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h0000000c, 1'b0, 32'hxxxxxxxx, 32'h00000008, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000008, 32'h00000008, 32'h0000000c, 5'h02, 32'h0000000c, 32'h00000004, 32'h00000008, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#789 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h01860186, 32'h0000000c, 32'hxxxxxxxx, 32'h00000008};
#790 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h00168000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h0000001d, 32'h0000001b, 32'h00000002, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001d, 32'h0000001b, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#790 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01860186, 32'h00000002, 32'hxxxxxxxx, 32'h0000001b};
#791 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ec, 32'h004a082a, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h00168000, 16'h0800, 1'b1, 5'b1x011, 1'b0, 32'h0000000c, 32'h00000010, 32'h00000001, 5'h01, 32'h00000001, 32'h0000082a, 32'h0000000c, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#791 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01860186, 32'h00000001, 32'hxxxxxxxx, 32'h00000010};
#792 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h0c6, 10'h000, 12'hfc6};
#792 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f0, 32'h1420fff9, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00168000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hfffffff9, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#792 bmem_addr <= 'h0206;
#792 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01860186, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#793 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h00000001, 32'h00168000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#793 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01860186, 32'h10010000, 32'h00000000, 32'h00000001};
#794 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h1001000c, 1'b0, 32'h00000023, 32'h0000000c, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h0000000c, 32'h1001000c, 5'h01, 32'h1001000c, 32'h00000821, 32'h10010000, 32'h0000000c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#794 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001b, 32'h01860186, 32'h1001000c, 32'h00000023, 32'h0000000c};
#795 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010014, 1'b0, 32'h0000001b, 32'h0000001d, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h1001000c, 32'h0000001d, 32'h10010014, 5'h08, 32'h0000001b, 32'h00000008, 32'h1001000c, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#795 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h0000001b, 32'h01860186, 32'h10010014, 32'h0000001b, 32'h0000001d};
#796 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000010, 1'b0, 32'hxxxxxxxx, 32'h0000000c, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h0000000c, 32'h0000000c, 32'h00000010, 5'h02, 32'h00000010, 32'h00000004, 32'h0000000c, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#796 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001b, 32'h01860186, 32'h00000010, 32'hxxxxxxxx, 32'h0000000c};
#796 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h0c7, 10'h000, 12'hfc6};
#796 bmem_addr <= 'h0207;
#797 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h00168000, 16'h0800, 1'b0, 5'b1xx01, 1'b1, 32'h0000001b, 32'h0000001b, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001b, 32'h0000001b, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#797 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001b, 32'h01860186, 32'h00000000, 32'hxxxxxxxx, 32'h0000001b};
#798 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f8, 32'h00021082, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h00168000, 16'h0800, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00000010, 32'h00000004, 5'h02, 32'h00000004, 32'h00001082, 32'h00000002, 32'h00000010, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#798 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001b, 32'h01860186, 32'h00000004, 32'hxxxxxxxx, 32'h00000010};
#799 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001fc, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h0040004c, 32'h0040004c, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'h1f, 32'h0040004c, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#799 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h0000001b, 32'h01860186, 32'h10010ffc, 32'h0040004c, 32'h0040004c};
#800 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01900190, 32'h10010ff8, 32'hxxxxxxxx, 32'h0000001b};
#800 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h0c8, 10'h000, 12'hfc6};
#800 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400200, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001b, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#800 bmem_addr <= 'h0208;
#801 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400204, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h0000001b, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001b, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#801 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01900190, 32'h10010ff4, 32'hxxxxxxxx, 32'h0000001b};
#802 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400208, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000010, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#802 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01900190, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000010};
#803 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040020c, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#803 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01900190, 32'h10011000, 32'h00000000, 32'h10010ff0};
#804 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400210, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00168000, 16'h0800, 1'b0, 5'bxxxxx, 1'bx, 32'h0040004c, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#804 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01900190, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#804 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h6, 10'h0c9, 10'h000, 12'hfc6};
#804 bmem_addr <= 'h0209;
#805 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h00028021, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000004, 32'h00000004, 5'h10, 32'h00000004, 32'hxxxx8021, 32'h00000000, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#805 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001c, 32'h01900190, 32'h00000004, 32'hxxxxxxxx, 32'h00000004};
#806 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h0c1000e2, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00168000, 16'h0800, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400054, 32'h000000e2, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#806 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01900190, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#807 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400388, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h1001000c, 32'h00168000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h1001000c, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#807 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01900190, 32'h10030000, 32'h0000001c, 32'h1001000c};
#808 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040038c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h00168000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#808 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01900190, 32'h10030000, 32'h0000001c, 32'h00000000};
#808 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hc, 4'h8, 10'h0ca, 10'h000, 12'hfc8};
#808 bmem_addr <= 'h020a;
#809 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400390, 32'hac200008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h00000000, 32'h00168000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#809 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001c, 32'h01900190, 32'h10030008, 32'hxxxxxxxx, 32'h00000000};
#810 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400394, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0800, 1'b0, 5'bxxxxx, 1'bx, 32'h00400054, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#810 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01900190, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#811 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400054, 32'h1200ffef, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h00000004, 32'h00000000, 32'h00000004, 5'hxx, 32'hxxxxxxxx, 32'hffffffef, 32'h00000004, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#811 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001c, 32'h01900190, 32'h00000004, 32'hxxxxxxxx, 32'h00000000};
#812 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'he, 4'hc, 10'h0cb, 10'h000, 12'hfec};
#812 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400058, 32'h20010001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h10030000, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h10030000, 32'h00000001, 5'h01, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#812 bmem_addr <= 'h020b;
#812 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01900190, 32'h00000001, 32'hxxxxxxxx, 32'h10030000};
#813 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040005c, 32'h14300005, 32'hfffffffd, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000004, 32'hfffffffd, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000001, 32'h00000004, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#813 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001c, 32'h01900190, 32'hfffffffd, 32'hxxxxxxxx, 32'h00000004};
#814 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400074, 32'h20010002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000001, 32'h00000002, 5'h01, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#814 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01900190, 32'h00000002, 32'hxxxxxxxx, 32'h00000001};
#815 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400078, 32'h14300005, 32'hfffffffe, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h00000002, 32'h00000004, 32'hfffffffe, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000002, 32'h00000004, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#815 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001c, 32'h01900190, 32'hfffffffe, 32'hxxxxxxxx, 32'h00000004};
#816 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0cc, 10'h000, 12'hfff};
#816 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400090, 32'h20010003, 32'h00000003, 1'b0, 32'hxxxxxxxx, 32'h00000002, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000002, 32'h00000003, 5'h01, 32'h00000003, 32'h00000003, 32'h00000000, 32'h00000003, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#816 bmem_addr <= 'h020c;
#816 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01900190, 32'h00000003, 32'hxxxxxxxx, 32'h00000002};
#817 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400094, 32'h14300005, 32'hffffffff, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h00000003, 32'h00000004, 32'hffffffff, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000003, 32'h00000004, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#817 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'h0040004c, 32'h0000001c, 32'h01900190, 32'hffffffff, 32'hxxxxxxxx, 32'h00000004};
#818 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000ac, 32'h20010004, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000003, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000003, 32'h00000004, 5'h01, 32'h00000004, 32'h00000004, 32'h00000000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#818 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001c, 32'h01900190, 32'h00000004, 32'hxxxxxxxx, 32'h00000003};
#819 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000b0, 32'h1430ffd8, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0800, 1'b0, 5'b1xx01, 1'b1, 32'h00000004, 32'h00000004, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'hffffffd8, 32'h00000004, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#819 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01900190, 32'h00000000, 32'hxxxxxxxx, 32'h00000004};
#820 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001c, 32'h019a019a, 32'h0000000f, 32'hxxxxxxxx, 32'h0000000e};
#820 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0cd, 10'h000, 12'hfff};
#820 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000b4, 32'h22520001, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h0000000e, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h0000000e, 32'h0000000e, 32'h0000000f, 5'h12, 32'h0000000f, 32'h00000001, 32'h0000000e, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#820 bmem_addr <= 'h020d;
#821 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000b8, 32'h2a41001e, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0800, 1'b1, 5'b1x011, 1'b0, 32'h0000000f, 32'h00000004, 32'h00000001, 5'h01, 32'h00000001, 32'h0000001e, 32'h0000000f, 32'h0000001e, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#821 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h019a019a, 32'h00000001, 32'hxxxxxxxx, 32'h00000004};
#822 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000bc, 32'h1420ffd5, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0800, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hffffffd5, 32'h00000001, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#822 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h019a019a, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#823 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h24040002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#823 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h019a019a, 32'h00000002, 32'hxxxxxxxx, 32'h0000000f};
#824 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00112821, 32'h00000016, 1'b0, 32'hxxxxxxxx, 32'h00000016, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000016, 32'h00000016, 5'h05, 32'h00000016, 32'h00002821, 32'h00000000, 32'h00000016, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#824 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h0000001c, 32'h019a019a, 32'h00000016, 32'hxxxxxxxx, 32'h00000016};
#824 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0ce, 10'h000, 12'hfff};
#824 bmem_addr <= 'h020e;
#825 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h00123021, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h0000000f, 5'h06, 32'h0000000f, 32'h00003021, 32'h00000000, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#825 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001c, 32'h019a019a, 32'h0000000f, 32'hxxxxxxxx, 32'h0000000f};
#826 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h0c10003e, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0800, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400024, 32'h0000003e, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#826 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h019a019a, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#827 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000f8, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#827 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h019a019a, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#828 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h0040004c, 32'h00400024, 32'h00000000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#828 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h0000001c, 32'h019a019a, 32'h10010ffc, 32'h0040004c, 32'h00400024};
#828 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'hf, 4'hf, 10'h0cf, 10'h000, 12'hfff};
#828 bmem_addr <= 'h020f;
#829 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h019a019a, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#829 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#830 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#830 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h019a019a, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#831 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#831 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h019a019a, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#832 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h0d0, 10'h000, 12'hccc};
#832 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'h00000001, 32'h00000000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000001, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#832 smem_addr <= 'h00d;
#832 bmem_addr <= 'h0300;
#832 charcode  <= 'h03;
#832 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h019a019a, 32'h10020000, 32'h00000000, 32'h00000001};
#833 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h0800, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'hxxxxxxxx, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#833 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h019a019a, 32'h10020000, 32'h00000000, 32'hxxxxxxxx};
#834 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h00064940, 32'h000001e0, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h000001e0, 5'h09, 32'h000001e0, 32'h00004940, 32'h00000005, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#834 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h019a019a, 32'h000001e0, 32'hxxxxxxxx, 32'h0000000f};
#835 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h000650c0, 32'h00000078, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000078, 5'h0a, 32'h00000078, 32'h000050c0, 32'h00000003, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#835 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h019a019a, 32'h00000078, 32'hxxxxxxxx, 32'h0000000f};
#836 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h0d1, 10'h000, 12'hccc};
#836 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h012a4820, 32'h00000258, 1'b0, 32'hxxxxxxxx, 32'h00000078, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h000001e0, 32'h00000078, 32'h00000258, 5'h09, 32'h00000258, 32'h00004820, 32'h000001e0, 32'h00000078, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#836 bmem_addr <= 'h0301;
#836 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h019a019a, 32'h00000258, 32'hxxxxxxxx, 32'h00000078};
#837 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h01254820, 32'h0000026e, 1'b0, 32'hxxxxxxxx, 32'h00000016, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000258, 32'h00000016, 32'h0000026e, 5'h09, 32'h0000026e, 32'h00004820, 32'h00000258, 32'h00000016, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#837 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h019a019a, 32'h0000026e, 32'hxxxxxxxx, 32'h00000016};
#838 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h00094880, 32'h000009b8, 1'b0, 32'hxxxxxxxx, 32'h0000026e, 32'h00000000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000026e, 32'h000009b8, 5'h09, 32'h000009b8, 32'h00004880, 32'h00000002, 32'h0000026e, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#838 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h019a019a, 32'h000009b8, 32'hxxxxxxxx, 32'h0000026e};
#839 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h01094020, 32'h100209b8, 1'b0, 32'h00000000, 32'h000009b8, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000009b8, 32'h100209b8, 5'h08, 32'h100209b8, 32'h00004020, 32'h10020000, 32'h000009b8, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#839 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h019a019a, 32'h100209b8, 32'h00000000, 32'h000009b8};
#840 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01a401a4, 32'h100209b8, 32'h00000000, 32'h00000002};
#840 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'had040000, 32'h100209b8, 1'b1, 32'h00000000, 32'h00000002, 32'h00000000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h100209b8, 32'h00000002, 32'h100209b8, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100209b8, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#840 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b1, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h0d2, 10'h000, 12'hccc};
#840 bmem_addr <= 'h0302;
#841 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001c, 32'h01a401a4, 32'h10010ffc, 32'h00400024, 32'h00400024};
#841 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h00400024, 32'h00400024, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'h1f, 32'h00400024, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#841 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h0d2, 10'h000, 12'hccc};
#842 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h100209b8, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100209b8, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#842 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01a401a4, 32'h10010ff8, 32'hxxxxxxxx, 32'h100209b8};
#843 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h000009b8, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000009b8, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#843 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01a401a4, 32'h10010ff4, 32'hxxxxxxxx, 32'h000009b8};
#844 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000078, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000078, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#844 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01a401a4, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000078};
#844 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hc, 4'hc, 4'hc, 10'h0d3, 10'h000, 12'hccc};
#844 bmem_addr <= 'h0303;
#845 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#845 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01a401a4, 32'h10011000, 32'h00000000, 32'h10010ff0};
#846 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400144, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0800, 1'b0, 5'bxxxxx, 1'bx, 32'h00400024, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#846 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01a401a4, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#847 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h0c1000d3, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0800, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400028, 32'h000000d3, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#847 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01a401a4, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#848 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040034c, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10020000, 32'h00000000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#848 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h0d4, 10'h000, 12'h999};
#848 bmem_addr <= 'h0304;
#848 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01a401a4, 32'h10030000, 32'h0000001c, 32'h10020000};
#849 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400350, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#849 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01a401a4, 32'h10030000, 32'h0000001c, 32'h00000000};
#850 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400354, 32'h8c220004, 32'h10030004, 1'b0, 32'h01a401a4, 32'h00000004, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000004, 32'h10030004, 5'h02, 32'h01a401a4, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#850 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001c, 32'h01a401a4, 32'h10030004, 32'h01a401a4, 32'h00000004};
#851 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400358, 32'h00021402, 32'h000001a4, 1'b0, 32'hxxxxxxxx, 32'h01a401a4, 32'h00000000, 16'h0800, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h01a401a4, 32'h000001a4, 5'h02, 32'h000001a4, 32'h00001402, 32'h00000010, 32'h01a401a4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#851 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01a401a4, 32'h000001a4, 32'hxxxxxxxx, 32'h01a401a4};
#852 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040035c, 32'h304201ff, 32'h000001a4, 1'b0, 32'hxxxxxxxx, 32'h000001a4, 32'h00000000, 16'h0800, 1'b1, 5'bx0000, 1'b0, 32'h000001a4, 32'h000001a4, 32'h000001a4, 5'h02, 32'h000001a4, 32'h000001ff, 32'h000001a4, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#852 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01a401a4, 32'h000001a4, 32'hxxxxxxxx, 32'h000001a4};
#852 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h0d5, 10'h000, 12'h999};
#852 bmem_addr <= 'h0305;
#853 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400360, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h0800, 1'b0, 5'bxxxxx, 1'bx, 32'h00400028, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#853 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01a401a4, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#854 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h00022300, 32'h001a4000, 1'b0, 32'h00000000, 32'h000001a4, 32'h00000000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000001a4, 32'h001a4000, 5'h04, 32'h001a4000, 32'h00002300, 32'h0000000c, 32'h000001a4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#854 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01a401a4, 32'h001a4000, 32'h00000000, 32'h000001a4};
#855 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h0c1000de, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h00000000, 16'h0800, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400030, 32'h000000de, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#855 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01a401a4, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#856 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400378, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10030000, 32'h00000000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#856 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'h9, 4'h9, 4'h9, 10'h0d6, 10'h000, 12'h999};
#856 bmem_addr <= 'h0306;
#856 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01a401a4, 32'h10030000, 32'h0000001c, 32'h10030000};
#857 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040037c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h00000000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#857 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01a401a4, 32'h10030000, 32'h0000001c, 32'h00000000};
#858 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400380, 32'hac240008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h001a4000, 32'h00000000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h001a4000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#858 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001c, 32'h01a401a4, 32'h10030008, 32'hxxxxxxxx, 32'h001a4000};
#859 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400384, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001a4000, 16'h0800, 1'b0, 5'bxxxxx, 1'bx, 32'h00400030, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#859 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01a401a4, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#860 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01ae01ae, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#860 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0d7, 10'h000, 12'hf20};
#860 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h0c1000d9, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h001a4000, 16'h0800, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400034, 32'h000000d9, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#860 bmem_addr <= 'h0307;
#861 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400364, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10030000, 32'h001a4000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#861 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ae01ae, 32'h10030000, 32'h0000001c, 32'h10030000};
#862 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400368, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h001a4000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#862 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ae01ae, 32'h10030000, 32'h0000001c, 32'h00000000};
#863 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040036c, 32'h8c220004, 32'h10030004, 1'b0, 32'h01ae01ae, 32'h000001a4, 32'h001a4000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h000001a4, 32'h10030004, 5'h02, 32'h01ae01ae, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#863 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001c, 32'h01ae01ae, 32'h10030004, 32'h01ae01ae, 32'h000001a4};
#864 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400370, 32'h304201ff, 32'h000001ae, 1'b0, 32'hxxxxxxxx, 32'h01ae01ae, 32'h001a4000, 16'h0800, 1'b1, 5'bx0000, 1'b0, 32'h01ae01ae, 32'h01ae01ae, 32'h000001ae, 5'h02, 32'h000001ae, 32'h000001ff, 32'h01ae01ae, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#864 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ae01ae, 32'h000001ae, 32'hxxxxxxxx, 32'h01ae01ae};
#864 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0d8, 10'h000, 12'hf20};
#864 bmem_addr <= 'h0308;
#865 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400374, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001a4000, 16'h0800, 1'b0, 5'bxxxxx, 1'bx, 32'h00400034, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#865 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01ae01ae, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#866 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h00021142, 32'h0000000d, 1'b0, 32'hxxxxxxxx, 32'h000001ae, 32'h001a4000, 16'h0800, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h000001ae, 32'h0000000d, 5'h02, 32'h0000000d, 32'h00001142, 32'h00000005, 32'h000001ae, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#866 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001c, 32'h01ae01ae, 32'h0000000d, 32'hxxxxxxxx, 32'h000001ae};
#867 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h24040001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h001a4000, 32'h001a4000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h001a4000, 32'h00000001, 5'h04, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#867 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ae01ae, 32'h00000001, 32'hxxxxxxxx, 32'h001a4000};
#868 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h00442004, 32'h00002000, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h001a4000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h0000000d, 32'h00000001, 32'h00002000, 5'h04, 32'h00002000, 32'h00002004, 32'h0000000d, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#868 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ae01ae, 32'h00002000, 32'hxxxxxxxx, 32'h00000001};
#868 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0d9, 10'h000, 12'hf20};
#868 bmem_addr <= 'h0309;
#869 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h0c1000e6, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h001a4000, 16'h0800, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h00400044, 32'h000000e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#869 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01ae01ae, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#870 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400398, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10030000, 32'h001a4000, 16'h0800, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#870 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ae01ae, 32'h10030000, 32'h0000001c, 32'h10030000};
#871 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040039c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h001a4000, 16'h0800, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#871 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ae01ae, 32'h10030000, 32'h0000001c, 32'h00000000};
#872 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0da, 10'h000, 12'hf20};
#872 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a0, 32'hac24000c, 32'h1003000c, 1'b1, 32'hxxxxxxxx, 32'h00002000, 32'h001a4000, 16'h0800, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00002000, 32'h1003000c, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10030000, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#872 bmem_addr <= 'h030a;
#872 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b1, 32'h00000003, 32'h00000023, 32'h0000001c, 32'h01ae01ae, 32'h1003000c, 32'hxxxxxxxx, 32'h00002000};
#873 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a4, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001a4000, 16'h2000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400044, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#873 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01ae01ae, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#874 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h2404000f, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h00002000, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00002000, 32'h0000000f, 5'h04, 32'h0000000f, 32'h0000000f, 32'h00000000, 32'h0000000f, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#874 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001c, 32'h01ae01ae, 32'h0000000f, 32'hxxxxxxxx, 32'h00002000};
#875 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h0c100066, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h001a4000, 16'h2000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000004, 32'hxxxxxxxx, 5'h1f, 32'h0040004c, 32'h00000066, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#875 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01ae01ae, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000004};
#876 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#876 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0db, 10'h000, 12'hf20};
#876 bmem_addr <= 'h030b;
#876 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01ae01ae, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#877 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h00400024, 32'h0040004c, 32'h001a4000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#877 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001c, 32'h01ae01ae, 32'h10010ffc, 32'h00400024, 32'h0040004c};
#877 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0db, 10'h000, 12'hf20};
#878 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01ae01ae, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#878 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h001a4000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#879 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h001a4000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#879 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01ae01ae, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#880 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01b801b8, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#880 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0dc, 10'h000, 12'hf20};
#880 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h001a4000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#880 bmem_addr <= 'h030c;
#881 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10030000, 32'h001a4000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#881 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01b801b8, 32'h10030000, 32'h0000001c, 32'h10030000};
#881 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0dc, 10'h000, 12'hf20};
#882 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#882 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01b801b8, 32'h10030000, 32'h0000001c, 32'h00000000};
#883 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8c220000, 32'h10030000, 1'b0, 32'h0000001c, 32'h0000000d, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h0000000d, 32'h10030000, 5'h02, 32'h0000001c, 32'h00000000, 32'h10030000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#883 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01b801b8, 32'h10030000, 32'h0000001c, 32'h0000000d};
#884 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h1040000f, 32'h0000001c, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001a4000, 16'h2000, 1'b0, 5'b1xx01, 1'b0, 32'h0000001c, 32'h00000000, 32'h0000001c, 5'hxx, 32'hxxxxxxxx, 32'h0000000f, 32'h0000001c, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#884 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000004b, 32'h0000001c, 32'h01b801b8, 32'h0000001c, 32'hxxxxxxxx, 32'h00000000};
#884 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0dd, 10'h000, 12'hf20};
#884 bmem_addr <= 'h030d;
#885 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h00024821, 32'h0000001c, 1'b0, 32'hxxxxxxxx, 32'h0000001c, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000001c, 32'h0000001c, 5'h09, 32'h0000001c, 32'h00004821, 32'h00000000, 32'h0000001c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#885 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000004b, 32'h0000001c, 32'h01b801b8, 32'h0000001c, 32'hxxxxxxxx, 32'h0000001c};
#886 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c0, 32'h24020000, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001c, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h0000001c, 32'h00000000, 5'h02, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#886 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01b801b8, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c};
#887 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c4, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10030000, 32'h001a4000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#887 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01b801b8, 32'h10010000, 32'h00000000, 32'h10030000};
#888 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c8, 32'h34280008, 32'h10010008, 1'b0, 32'h0000001c, 32'hxxxxxxxx, 32'h001a4000, 16'h2000, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010008, 5'h08, 32'h10010008, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#888 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001c, 32'h01b801b8, 32'h10010008, 32'h0000001c, 32'hxxxxxxxx};
#888 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0de, 10'h000, 12'hf20};
#888 bmem_addr <= 'h030e;
#889 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001cc, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h001a4000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#889 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01b801b8, 32'h10010000, 32'h00000000, 32'h10010000};
#890 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d0, 32'h342a0018, 32'h10010018, 1'b0, 32'h0000003b, 32'hxxxxxxxx, 32'h001a4000, 16'h2000, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010018, 5'h0a, 32'h10010018, 32'h00000018, 32'h10010000, 32'h00000018, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#890 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h0000001c, 32'h01b801b8, 32'h10010018, 32'h0000003b, 32'hxxxxxxxx};
#891 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d4, 32'h01485022, 32'h00000010, 1'b0, 32'hxxxxxxxx, 32'h10010008, 32'h001a4000, 16'h2000, 1'b1, 5'b1xx01, 1'b0, 32'h10010018, 32'h10010008, 32'h00000010, 5'h0a, 32'h00000010, 32'h00005022, 32'h10010018, 32'h10010008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#891 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001c, 32'h01b801b8, 32'h00000010, 32'hxxxxxxxx, 32'h10010008};
#892 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h001a4000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#892 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01b801b8, 32'h10010000, 32'h00000000, 32'h10010000};
#892 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0df, 10'h000, 12'hf20};
#892 bmem_addr <= 'h030f;
#893 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#893 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01b801b8, 32'h10010000, 32'h00000000, 32'h00000000};
#894 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010008, 1'b0, 32'h0000001c, 32'h10010008, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h10010008, 32'h10010008, 5'h08, 32'h0000001c, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#894 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001c, 32'h01b801b8, 32'h10010008, 32'h0000001c, 32'h10010008};
#895 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000004, 5'h02, 32'h00000004, 32'h00000004, 32'h00000000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#895 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001c, 32'h01b801b8, 32'h00000004, 32'hxxxxxxxx, 32'h00000000};
#896 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001c, 32'h001a4000, 16'h2000, 1'b0, 5'b1xx01, 1'b1, 32'h0000001c, 32'h0000001c, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001c, 32'h0000001c, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#896 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01b801b8, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c};
#896 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e0, 10'h000, 12'hf20};
#896 smem_addr <= 'h00e;
#896 bmem_addr <= 'h0000;
#896 charcode  <= 'h00;
#897 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f8, 32'h00021082, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h001a4000, 16'h2000, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00000004, 32'h00000001, 5'h02, 32'h00000001, 32'h00001082, 32'h00000002, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#897 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01b801b8, 32'h00000001, 32'hxxxxxxxx, 32'h00000004};
#898 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001fc, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h0040004c, 32'h0040004c, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'h1f, 32'h0040004c, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#898 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h0000001c, 32'h01b801b8, 32'h10010ffc, 32'h0040004c, 32'h0040004c};
#899 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400200, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h0000001c, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001c, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#899 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01b801b8, 32'h10010ff8, 32'hxxxxxxxx, 32'h0000001c};
#900 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01c201c2, 32'h10010ff4, 32'hxxxxxxxx, 32'h0000001c};
#900 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400204, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h0000001c, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001c, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#900 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e1, 10'h000, 12'hf20};
#900 bmem_addr <= 'h0001;
#901 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400208, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000010, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#901 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01c201c2, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000010};
#902 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040020c, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#902 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01c201c2, 32'h10011000, 32'h00000000, 32'h10010ff0};
#903 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400210, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001a4000, 16'h2000, 1'b0, 5'bxxxxx, 1'bx, 32'h0040004c, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#903 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01c201c2, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#904 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e2, 10'h000, 12'hf20};
#904 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h00028021, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000001, 32'h00000001, 5'h10, 32'h00000001, 32'hxxxx8021, 32'h00000000, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#904 bmem_addr <= 'h0002;
#904 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01c201c2, 32'h00000001, 32'hxxxxxxxx, 32'h00000001};
#905 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h0c1000e2, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h001a4000, 16'h2000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000001, 32'hxxxxxxxx, 5'h1f, 32'h00400054, 32'h000000e2, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#905 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01c201c2, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000001};
#906 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400388, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10010000, 32'h001a4000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#906 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01c201c2, 32'h10030000, 32'h0000001c, 32'h10010000};
#907 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040038c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h001a4000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#907 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01c201c2, 32'h10030000, 32'h0000001c, 32'h00000000};
#908 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e3, 10'h000, 12'hf20};
#908 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400390, 32'hac200008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h00000000, 32'h001a4000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#908 bmem_addr <= 'h0003;
#908 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001c, 32'h01c201c2, 32'h10030008, 32'hxxxxxxxx, 32'h00000000};
#909 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400394, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h2000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400054, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#909 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01c201c2, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#910 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400054, 32'h1200ffef, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h2000, 1'b0, 5'b1xx01, 1'b0, 32'h00000001, 32'h00000000, 32'h00000001, 5'hxx, 32'hxxxxxxxx, 32'hffffffef, 32'h00000001, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#910 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01c201c2, 32'h00000001, 32'hxxxxxxxx, 32'h00000000};
#911 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400058, 32'h20010001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h10030000, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h10030000, 32'h00000001, 5'h01, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#911 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01c201c2, 32'h00000001, 32'hxxxxxxxx, 32'h10030000};
#912 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040005c, 32'h14300005, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00000000, 16'h2000, 1'b0, 5'b1xx01, 1'b1, 32'h00000001, 32'h00000001, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000005, 32'h00000001, 32'h00000001, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#912 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01c201c2, 32'h00000000, 32'hxxxxxxxx, 32'h00000001};
#912 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e4, 10'h000, 12'hf20};
#912 bmem_addr <= 'h0004;
#913 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400060, 32'h2231ffff, 32'h00000015, 1'b0, 32'hxxxxxxxx, 32'h00000016, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h00000016, 32'h00000016, 32'h00000015, 5'h11, 32'h00000015, 32'hffffffff, 32'h00000016, 32'hffffffff, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#913 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h0000001c, 32'h01c201c2, 32'h00000015, 32'hxxxxxxxx, 32'h00000016};
#914 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400064, 32'h0220082a, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h2000, 1'b1, 5'b1x011, 1'b1, 32'h00000015, 32'h00000000, 32'h00000000, 5'h01, 32'h00000000, 32'h0000082a, 32'h00000015, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#914 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01c201c2, 32'h00000000, 32'hxxxxxxxx, 32'h00000000};
#915 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400068, 32'h1020ffea, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h2000, 1'b0, 5'b1xx01, 1'b1, 32'h00000000, 32'h00000000, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'hffffffea, 32'h00000000, 32'h00000000, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#916 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e5, 10'h000, 12'hf20};
#916 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400014, 32'h24040002, 32'h00000002, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000002, 5'h04, 32'h00000002, 32'h00000002, 32'h00000000, 32'h00000002, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#916 bmem_addr <= 'h0005;
#916 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01c201c2, 32'h00000002, 32'hxxxxxxxx, 32'h0000000f};
#917 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400018, 32'h00112821, 32'h00000015, 1'b0, 32'hxxxxxxxx, 32'h00000015, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000015, 32'h00000015, 5'h05, 32'h00000015, 32'h00002821, 32'h00000000, 32'h00000015, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#917 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001b, 32'h0000001c, 32'h01c201c2, 32'h00000015, 32'hxxxxxxxx, 32'h00000015};
#918 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040001c, 32'h00123021, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000000f, 32'h0000000f, 5'h06, 32'h0000000f, 32'h00003021, 32'h00000000, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#918 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001c, 32'h01c201c2, 32'h0000000f, 32'hxxxxxxxx, 32'h0000000f};
#919 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400020, 32'h0c10003e, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00000000, 16'h2000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000001, 32'hxxxxxxxx, 5'h1f, 32'h00400024, 32'h0000003e, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#919 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01c201c2, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000001};
#920 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01cc01cc, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#920 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000f8, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#920 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e6, 10'h000, 12'hf20};
#920 bmem_addr <= 'h0006;
#921 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004000fc, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h0040004c, 32'h00400024, 32'h00000000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#921 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h0000001c, 32'h01cc01cc, 32'h10010ffc, 32'h0040004c, 32'h00400024};
#921 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e6, 10'h000, 12'hf20};
#922 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01cc01cc, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#922 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400100, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#923 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400104, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#923 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01cc01cc, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#924 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e7, 10'h000, 12'hf20};
#924 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400108, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#924 bmem_addr <= 'h0007;
#924 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01cc01cc, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#925 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040010c, 32'h3c011002, 32'h10020000, 1'b0, 32'h00000000, 32'h00000000, 32'h00000000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h00000000, 32'h10020000, 5'h01, 32'h10020000, 32'h00001002, 32'h00000010, 32'h00001002, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#925 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01cc01cc, 32'h10020000, 32'h00000000, 32'h00000000};
#925 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e7, 10'h000, 12'hf20};
#926 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400110, 32'h34280000, 32'h10020000, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h00000000, 16'h2000, 1'b1, 5'bx0100, 1'b0, 32'h10020000, 32'hxxxxxxxx, 32'h10020000, 5'h08, 32'h10020000, 32'h00000000, 32'h10020000, 32'h00000000, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#926 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01cc01cc, 32'h10020000, 32'h00000000, 32'hxxxxxxxx};
#927 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400114, 32'h00064940, 32'h000001e0, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h000001e0, 5'h09, 32'h000001e0, 32'h00004940, 32'h00000005, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#927 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01cc01cc, 32'h000001e0, 32'hxxxxxxxx, 32'h0000000f};
#928 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e8, 10'h000, 12'hf20};
#928 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400118, 32'h000650c0, 32'h00000078, 1'b0, 32'hxxxxxxxx, 32'h0000000f, 32'h00000000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000000f, 32'h00000078, 5'h0a, 32'h00000078, 32'h000050c0, 32'h00000003, 32'h0000000f, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#928 bmem_addr <= 'h0008;
#928 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01cc01cc, 32'h00000078, 32'hxxxxxxxx, 32'h0000000f};
#929 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040011c, 32'h012a4820, 32'h00000258, 1'b0, 32'hxxxxxxxx, 32'h00000078, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h000001e0, 32'h00000078, 32'h00000258, 5'h09, 32'h00000258, 32'h00004820, 32'h000001e0, 32'h00000078, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#929 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01cc01cc, 32'h00000258, 32'hxxxxxxxx, 32'h00000078};
#930 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400120, 32'h01254820, 32'h0000026d, 1'b0, 32'hxxxxxxxx, 32'h00000015, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h00000258, 32'h00000015, 32'h0000026d, 5'h09, 32'h0000026d, 32'h00004820, 32'h00000258, 32'h00000015, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#930 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01cc01cc, 32'h0000026d, 32'hxxxxxxxx, 32'h00000015};
#931 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400124, 32'h00094880, 32'h000009b4, 1'b0, 32'hxxxxxxxx, 32'h0000026d, 32'h00000000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h0000026d, 32'h000009b4, 5'h09, 32'h000009b4, 32'h00004880, 32'h00000002, 32'h0000026d, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#931 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000000, 32'h0000001c, 32'h01cc01cc, 32'h000009b4, 32'hxxxxxxxx, 32'h0000026d};
#932 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400128, 32'h01094020, 32'h100209b4, 1'b0, 32'h00000003, 32'h000009b4, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10020000, 32'h000009b4, 32'h100209b4, 5'h08, 32'h100209b4, 32'h00004020, 32'h10020000, 32'h000009b4, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#932 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000000, 32'h0000001c, 32'h01cc01cc, 32'h100209b4, 32'h00000003, 32'h000009b4};
#932 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e9, 10'h000, 12'hf20};
#932 bmem_addr <= 'h0009;
#933 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040012c, 32'had040000, 32'h100209b4, 1'b1, 32'h00000003, 32'h00000002, 32'h00000000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h100209b4, 32'h00000002, 32'h100209b4, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h100209b4, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#933 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000000, 32'h0000001c, 32'h01cc01cc, 32'h100209b4, 32'h00000003, 32'h00000002};
#933 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b1, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e9, 10'h000, 12'hf20};
#934 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001c, 32'h01cc01cc, 32'h10010ffc, 32'h00400024, 32'h00400024};
#934 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400130, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h00400024, 32'h00400024, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00400024, 32'h10010ffc, 5'h1f, 32'h00400024, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#934 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0e9, 10'h000, 12'hf20};
#935 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400134, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h100209b4, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h100209b4, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#935 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01cc01cc, 32'h10010ff8, 32'hxxxxxxxx, 32'h100209b4};
#936 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400138, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h000009b4, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h000009b4, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#936 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01cc01cc, 32'h10010ff4, 32'hxxxxxxxx, 32'h000009b4};
#936 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0ea, 10'h000, 12'hf20};
#936 bmem_addr <= 'h000a;
#937 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040013c, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000078, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000078, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#937 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01cc01cc, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000078};
#938 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400140, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#938 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01cc01cc, 32'h10011000, 32'h00000000, 32'h10010ff0};
#939 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400144, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h2000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400024, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#939 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01cc01cc, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#940 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01d601d6, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000001};
#940 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0eb, 10'h000, 12'hf20};
#940 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400024, 32'h0c1000d3, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00000000, 16'h2000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000001, 32'hxxxxxxxx, 5'h1f, 32'h00400028, 32'h000000d3, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#940 bmem_addr <= 'h000b;
#941 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040034c, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10020000, 32'h00000000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10020000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#941 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01d601d6, 32'h10030000, 32'h0000001c, 32'h10020000};
#942 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400350, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#942 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01d601d6, 32'h10030000, 32'h0000001c, 32'h00000000};
#943 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400354, 32'h8c220004, 32'h10030004, 1'b0, 32'h01d601d6, 32'h00000001, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000001, 32'h10030004, 5'h02, 32'h01d601d6, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#943 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001c, 32'h01d601d6, 32'h10030004, 32'h01d601d6, 32'h00000001};
#944 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400358, 32'h00021402, 32'h000001d6, 1'b0, 32'hxxxxxxxx, 32'h01d601d6, 32'h00000000, 16'h2000, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h01d601d6, 32'h000001d6, 5'h02, 32'h000001d6, 32'h00001402, 32'h00000010, 32'h01d601d6, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#944 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01d601d6, 32'h000001d6, 32'hxxxxxxxx, 32'h01d601d6};
#944 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0ec, 10'h000, 12'hf20};
#944 bmem_addr <= 'h000c;
#945 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040035c, 32'h304201ff, 32'h000001d6, 1'b0, 32'hxxxxxxxx, 32'h000001d6, 32'h00000000, 16'h2000, 1'b1, 5'bx0000, 1'b0, 32'h000001d6, 32'h000001d6, 32'h000001d6, 5'h02, 32'h000001d6, 32'h000001ff, 32'h000001d6, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#945 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01d601d6, 32'h000001d6, 32'hxxxxxxxx, 32'h000001d6};
#946 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400360, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h00000000, 16'h2000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400028, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#946 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01d601d6, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#947 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400028, 32'h00022300, 32'h001d6000, 1'b0, 32'h00000000, 32'h000001d6, 32'h00000000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h000001d6, 32'h001d6000, 5'h04, 32'h001d6000, 32'h00002300, 32'h0000000c, 32'h000001d6, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#947 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01d601d6, 32'h001d6000, 32'h00000000, 32'h000001d6};
#948 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0ed, 10'h000, 12'hf20};
#948 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040002c, 32'h0c1000de, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h00000000, 16'h2000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000001, 32'hxxxxxxxx, 5'h1f, 32'h00400030, 32'h000000de, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#948 bmem_addr <= 'h000d;
#948 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01d601d6, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000001};
#949 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400378, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10030000, 32'h00000000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#949 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01d601d6, 32'h10030000, 32'h0000001c, 32'h10030000};
#950 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040037c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h00000000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#950 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01d601d6, 32'h10030000, 32'h0000001c, 32'h00000000};
#951 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400380, 32'hac240008, 32'h10030008, 1'b1, 32'hxxxxxxxx, 32'h001d6000, 32'h00000000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h001d6000, 32'h10030008, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10030000, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#951 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b1, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001c, 32'h01d601d6, 32'h10030008, 32'hxxxxxxxx, 32'h001d6000};
#952 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400384, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001d6000, 16'h2000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400030, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#952 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0ee, 10'h000, 12'hf20};
#952 bmem_addr <= 'h000e;
#952 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01d601d6, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#953 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400030, 32'h0c1000d9, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h001d6000, 16'h2000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000001, 32'hxxxxxxxx, 5'h1f, 32'h00400034, 32'h000000d9, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#953 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01d601d6, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000001};
#954 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400364, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10030000, 32'h001d6000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#954 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01d601d6, 32'h10030000, 32'h0000001c, 32'h10030000};
#955 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400368, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h001d6000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#955 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01d601d6, 32'h10030000, 32'h0000001c, 32'h00000000};
#956 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0ef, 10'h000, 12'hf20};
#956 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040036c, 32'h8c220004, 32'h10030004, 1'b0, 32'h01d601d6, 32'h000001d6, 32'h001d6000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h000001d6, 32'h10030004, 5'h02, 32'h01d601d6, 32'h00000004, 32'h10030000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#956 bmem_addr <= 'h000f;
#956 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001c, 32'h01d601d6, 32'h10030004, 32'h01d601d6, 32'h000001d6};
#957 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400370, 32'h304201ff, 32'h000001d6, 1'b0, 32'hxxxxxxxx, 32'h01d601d6, 32'h001d6000, 16'h2000, 1'b1, 5'bx0000, 1'b0, 32'h01d601d6, 32'h01d601d6, 32'h000001d6, 5'h02, 32'h000001d6, 32'h000001ff, 32'h01d601d6, 32'h000001ff, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#957 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01d601d6, 32'h000001d6, 32'hxxxxxxxx, 32'h01d601d6};
#958 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400374, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001d6000, 16'h2000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400034, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#958 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01d601d6, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#959 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400034, 32'h00021142, 32'h0000000e, 1'b0, 32'hxxxxxxxx, 32'h000001d6, 32'h001d6000, 16'h2000, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h000001d6, 32'h0000000e, 5'h02, 32'h0000000e, 32'h00001142, 32'h00000005, 32'h000001d6, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#959 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001c, 32'h01d601d6, 32'h0000000e, 32'hxxxxxxxx, 32'h000001d6};
#960 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01e001e0, 32'h00000001, 32'hxxxxxxxx, 32'h001d6000};
#960 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400038, 32'h24040001, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h001d6000, 32'h001d6000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h001d6000, 32'h00000001, 5'h04, 32'h00000001, 32'h00000001, 32'h00000000, 32'h00000001, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#960 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f0, 10'h000, 12'hf20};
#960 smem_addr <= 'h00f;
#960 bmem_addr <= 'h0000;
#961 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040003c, 32'h00442004, 32'h00004000, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h001d6000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h0000000e, 32'h00000001, 32'h00004000, 5'h04, 32'h00004000, 32'h00002004, 32'h0000000e, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#961 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01e001e0, 32'h00004000, 32'hxxxxxxxx, 32'h00000001};
#962 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400040, 32'h0c1000e6, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h001d6000, 16'h2000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000001, 32'hxxxxxxxx, 5'h1f, 32'h00400044, 32'h000000e6, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#962 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01e001e0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000001};
#963 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400398, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10030000, 32'h001d6000, 16'h2000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#963 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01e001e0, 32'h10030000, 32'h0000001c, 32'h10030000};
#964 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f1, 10'h000, 12'hf20};
#964 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040039c, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h001d6000, 16'h2000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#964 bmem_addr <= 'h0001;
#964 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01e001e0, 32'h10030000, 32'h0000001c, 32'h00000000};
#965 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a0, 32'hac24000c, 32'h1003000c, 1'b1, 32'hxxxxxxxx, 32'h00004000, 32'h001d6000, 16'h2000, 1'b0, 5'b0xx01, 1'b0, 32'h10030000, 32'h00004000, 32'h1003000c, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10030000, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#965 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b1, 32'h00000003, 32'h00000023, 32'h0000001c, 32'h01e001e0, 32'h1003000c, 32'hxxxxxxxx, 32'h00004000};
#966 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004003a4, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001d6000, 16'h4000, 1'b0, 5'bxxxxx, 1'bx, 32'h00400044, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#966 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01e001e0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#967 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400044, 32'h2404000f, 32'h0000000f, 1'b0, 32'hxxxxxxxx, 32'h00004000, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00004000, 32'h0000000f, 5'h04, 32'h0000000f, 32'h0000000f, 32'h00000000, 32'h0000000f, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#967 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000003, 32'h00000023, 32'h0000001c, 32'h01e001e0, 32'h0000000f, 32'hxxxxxxxx, 32'h00004000};
#968 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400048, 32'h0c100066, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h001d6000, 16'h4000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000001, 32'hxxxxxxxx, 5'h1f, 32'h0040004c, 32'h00000066, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#968 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01e001e0, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000001};
#968 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f2, 10'h000, 12'hf20};
#968 bmem_addr <= 'h0002;
#969 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400198, 32'h23bdfff0, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h10011000, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h10011000, 32'h10011000, 32'h10010ff0, 5'h1d, 32'h10010ff0, 32'hfffffff0, 32'h10011000, 32'hfffffff0, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#969 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01e001e0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10011000};
#970 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040019c, 32'hafbf000c, 32'h10010ffc, 1'b1, 32'h00400024, 32'h0040004c, 32'h001d6000, 16'h4000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'hxx, 32'hxxxxxxxx, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#970 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00400024, 32'h0000001c, 32'h01e001e0, 32'h10010ffc, 32'h00400024, 32'h0040004c};
#970 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f2, 10'h000, 12'hf20};
#971 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01e001e0, 32'h10010ff8, 32'hxxxxxxxx, 32'hxxxxxxxx};
#971 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a0, 32'hafa80008, 32'h10010ff8, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h001d6000, 16'h4000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff8, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#972 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b1, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f3, 10'h000, 12'hf20};
#972 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a4, 32'hafa90004, 32'h10010ff4, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h001d6000, 16'h4000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff4, 5'hxx, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#972 bmem_addr <= 'h0003;
#972 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01e001e0, 32'h10010ff4, 32'hxxxxxxxx, 32'hxxxxxxxx};
#973 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001a8, 32'hafaa0000, 32'h10010ff0, 1'b1, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h001d6000, 16'h4000, 1'b0, 5'b0xx01, 1'b0, 32'h10010ff0, 32'hxxxxxxxx, 32'h10010ff0, 5'hxx, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b1, 2'bxx, 1'b1, 2'b00};
#973 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01e001e0, 32'h10010ff0, 32'hxxxxxxxx, 32'hxxxxxxxx};
#974 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001ac, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10030000, 32'h001d6000, 16'h4000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#974 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01e001e0, 32'h10030000, 32'h0000001c, 32'h10030000};
#974 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f3, 10'h000, 12'hf20};
#975 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b0, 32'h00200821, 32'h10030000, 1'b0, 32'h0000001c, 32'h00000000, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h00000000, 32'h10030000, 5'h01, 32'h10030000, 32'h00000821, 32'h10030000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#975 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01e001e0, 32'h10030000, 32'h0000001c, 32'h00000000};
#976 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f4, 10'h000, 12'hf20};
#976 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b4, 32'h8c220000, 32'h10030000, 1'b0, 32'h0000001c, 32'h0000000e, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h10030000, 32'h0000000e, 32'h10030000, 5'h02, 32'h0000001c, 32'h00000000, 32'h10030000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#976 bmem_addr <= 'h0004;
#976 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01e001e0, 32'h10030000, 32'h0000001c, 32'h0000000e};
#977 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001b8, 32'h1040000f, 32'h0000001c, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001d6000, 16'h4000, 1'b0, 5'b1xx01, 1'b0, 32'h0000001c, 32'h00000000, 32'h0000001c, 5'hxx, 32'hxxxxxxxx, 32'h0000000f, 32'h0000001c, 32'h00000000, 2'b00, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#977 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000004b, 32'h0000001c, 32'h01e001e0, 32'h0000001c, 32'hxxxxxxxx, 32'h00000000};
#978 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001bc, 32'h00024821, 32'h0000001c, 1'b0, 32'hxxxxxxxx, 32'h0000001c, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h0000001c, 32'h0000001c, 5'h09, 32'h0000001c, 32'h00004821, 32'h00000000, 32'h0000001c, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#978 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000004b, 32'h0000001c, 32'h01e001e0, 32'h0000001c, 32'hxxxxxxxx, 32'h0000001c};
#979 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c0, 32'h24020000, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001c, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b1, 32'h00000000, 32'h0000001c, 32'h00000000, 5'h02, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#979 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01e001e0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c};
#980 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ea01ea, 32'h10010000, 32'h00000000, 32'h10030000};
#980 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c4, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10030000, 32'h001d6000, 16'h4000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10030000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#980 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f5, 10'h000, 12'hf20};
#980 bmem_addr <= 'h0005;
#981 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001c8, 32'h34280008, 32'h10010008, 1'b0, 32'h0000001c, 32'hxxxxxxxx, 32'h001d6000, 16'h4000, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010008, 5'h08, 32'h10010008, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#981 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001c, 32'h01ea01ea, 32'h10010008, 32'h0000001c, 32'hxxxxxxxx};
#982 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001cc, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h001d6000, 16'h4000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#982 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ea01ea, 32'h10010000, 32'h00000000, 32'h10010000};
#983 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d0, 32'h342a0018, 32'h10010018, 1'b0, 32'h0000003b, 32'hxxxxxxxx, 32'h001d6000, 16'h4000, 1'b1, 5'bx0100, 1'b0, 32'h10010000, 32'hxxxxxxxx, 32'h10010018, 5'h0a, 32'h10010018, 32'h00000018, 32'h10010000, 32'h00000018, 2'b00, 2'b01, 1'b0, 1'b1, 2'b01, 1'b0, 2'b00};
#983 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h0000003b, 32'h0000001c, 32'h01ea01ea, 32'h10010018, 32'h0000003b, 32'hxxxxxxxx};
#984 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d4, 32'h01485022, 32'h00000010, 1'b0, 32'hxxxxxxxx, 32'h10010008, 32'h001d6000, 16'h4000, 1'b1, 5'b1xx01, 1'b0, 32'h10010018, 32'h10010008, 32'h00000010, 5'h0a, 32'h00000010, 32'h00005022, 32'h10010018, 32'h10010008, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#984 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0000001d, 32'h0000001c, 32'h01ea01ea, 32'h00000010, 32'hxxxxxxxx, 32'h10010008};
#984 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f6, 10'h000, 12'hf20};
#984 bmem_addr <= 'h0006;
#985 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001d8, 32'h3c011001, 32'h10010000, 1'b0, 32'h00000000, 32'h10010000, 32'h001d6000, 16'h4000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10010000, 5'h01, 32'h10010000, 32'h00001001, 32'h00000010, 32'h00001001, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#985 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ea01ea, 32'h10010000, 32'h00000000, 32'h10010000};
#986 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001dc, 32'h00220821, 32'h10010000, 1'b0, 32'h00000000, 32'h00000000, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h00000000, 32'h10010000, 5'h01, 32'h10010000, 32'h00000821, 32'h10010000, 32'h00000000, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#986 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ea01ea, 32'h10010000, 32'h00000000, 32'h00000000};
#987 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e0, 32'h8c280008, 32'h10010008, 1'b0, 32'h0000001c, 32'h10010008, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h10010000, 32'h10010008, 32'h10010008, 5'h08, 32'h0000001c, 32'h00000008, 32'h10010000, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#987 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000002, 32'h0000001c, 32'h0000001c, 32'h01ea01ea, 32'h10010008, 32'h0000001c, 32'h10010008};
#988 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e4, 32'h20420004, 32'h00000004, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000000, 32'h00000004, 5'h02, 32'h00000004, 32'h00000004, 32'h00000000, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#988 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000001, 32'h00000003, 32'h0000001c, 32'h01ea01ea, 32'h00000004, 32'hxxxxxxxx, 32'h00000000};
#988 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f7, 10'h000, 12'hf20};
#988 bmem_addr <= 'h0007;
#989 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001e8, 32'h11090003, 32'h00000000, 1'b0, 32'hxxxxxxxx, 32'h0000001c, 32'h001d6000, 16'h4000, 1'b0, 5'b1xx01, 1'b1, 32'h0000001c, 32'h0000001c, 32'h00000000, 5'hxx, 32'hxxxxxxxx, 32'h00000003, 32'h0000001c, 32'h0000001c, 2'b01, 2'bxx, 1'b1, 1'b0, 2'bxx, 1'b0, 2'b00};
#989 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ea01ea, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c};
#990 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001f8, 32'h00021082, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000004, 32'h001d6000, 16'h4000, 1'b1, 5'bx1010, 1'b0, 32'h00000000, 32'h00000004, 32'h00000001, 5'h02, 32'h00000001, 32'h00001082, 32'h00000002, 32'h00000004, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b01};
#990 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ea01ea, 32'h00000001, 32'hxxxxxxxx, 32'h00000004};
#991 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h004001fc, 32'h8fbf000c, 32'h10010ffc, 1'b0, 32'h0040004c, 32'h0040004c, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0040004c, 32'h10010ffc, 5'h1f, 32'h0040004c, 32'h0000000c, 32'h10010ff0, 32'h0000000c, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#991 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h0040004c, 32'h0000001c, 32'h01ea01ea, 32'h10010ffc, 32'h0040004c, 32'h0040004c};
#992 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f8, 10'h000, 12'hf20};
#992 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400200, 32'h8fa80008, 32'h10010ff8, 1'b0, 32'hxxxxxxxx, 32'h0000001c, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001c, 32'h10010ff8, 5'h08, 32'hxxxxxxxx, 32'h00000008, 32'h10010ff0, 32'h00000008, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#992 bmem_addr <= 'h0008;
#992 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01ea01ea, 32'h10010ff8, 32'hxxxxxxxx, 32'h0000001c};
#993 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400204, 32'h8fa90004, 32'h10010ff4, 1'b0, 32'hxxxxxxxx, 32'h0000001c, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h0000001c, 32'h10010ff4, 5'h09, 32'hxxxxxxxx, 32'h00000004, 32'h10010ff0, 32'h00000004, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#993 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01ea01ea, 32'h10010ff4, 32'hxxxxxxxx, 32'h0000001c};
#994 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400208, 32'h8faa0000, 32'h10010ff0, 1'b0, 32'hxxxxxxxx, 32'h00000010, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h00000010, 32'h10010ff0, 5'h0a, 32'hxxxxxxxx, 32'h00000000, 32'h10010ff0, 32'h00000000, 2'b00, 2'b01, 1'b1, 1'b1, 2'b10, 1'b0, 2'b00};
#994 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'hxxxxxxxx, 32'h0000001c, 32'h01ea01ea, 32'h10010ff0, 32'hxxxxxxxx, 32'h00000010};
#995 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040020c, 32'h23bd0010, 32'h10011000, 1'b0, 32'h00000000, 32'h10010ff0, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h10010ff0, 32'h10010ff0, 32'h10011000, 5'h1d, 32'h10011000, 32'h00000010, 32'h10010ff0, 32'h00000010, 2'b00, 2'b01, 1'b1, 1'b1, 2'b01, 1'b0, 2'b00};
#995 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ea01ea, 32'h10011000, 32'h00000000, 32'h10010ff0};
#996 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400210, 32'h03e00008, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000000, 32'h001d6000, 16'h4000, 1'b0, 5'bxxxxx, 1'bx, 32'h0040004c, 32'h00000000, 32'hxxxxxxxx, 5'hxx, 32'hxxxxxxxx, 32'h00000008, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b11, 2'bxx, 1'bx, 1'bx, 2'bxx, 1'b0, 2'bxx};
#996 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01ea01ea, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000000};
#996 {dmem_wr, smem_wr, hsync, vsync, red, green, blue, x, y, bmem_color} <= {1'b0, 1'b0, 1'b1, 1'b1, 4'hf, 4'h2, 4'h0, 10'h0f9, 10'h000, 12'hf20};
#996 bmem_addr <= 'h0009;
#997 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h0040004c, 32'h00028021, 32'h00000001, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h001d6000, 16'h4000, 1'b1, 5'b0xx01, 1'b0, 32'h00000000, 32'h00000001, 32'h00000001, 5'h10, 32'h00000001, 32'hxxxx8021, 32'h00000000, 32'h00000001, 2'b00, 2'b00, 1'bx, 1'b0, 2'b01, 1'b0, 2'b00};
#997 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ea01ea, 32'h00000001, 32'hxxxxxxxx, 32'h00000001};
#998 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400050, 32'h0c1000e2, 32'hxxxxxxxx, 1'b0, 32'hxxxxxxxx, 32'h00000001, 32'h001d6000, 16'h4000, 1'b1, 5'bxxxxx, 1'bx, 32'h00000000, 32'h00000001, 32'hxxxxxxxx, 5'h1f, 32'h00400054, 32'h000000e2, 32'hxxxxxxxx, 32'hxxxxxxxx, 2'b10, 2'b10, 1'bx, 1'bx, 2'b00, 1'b0, 2'bxx};
#998 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h000000Xx, 32'hxxxxxxxx, 32'h0000001c, 32'h01ea01ea, 32'hxxxxxxxx, 32'hxxxxxxxx, 32'h00000001};
#999 {pc, instr, mem_addr, mem_wr, mem_readdata, mem_writedata, period, LED, werf, alufn, Z, ReadData1, ReadData2, alu_result, reg_writeaddr, reg_writedata, signImm, aluA, aluB, pcsel, wasel, sgnext, bsel, wdsel, wr, asel} <= {32'h00400388, 32'h3c011003, 32'h10030000, 1'b0, 32'h0000001c, 32'h10010000, 32'h001d6000, 16'h4000, 1'b1, 5'bx0010, 1'b0, 32'h00000000, 32'h10010000, 32'h10030000, 5'h01, 32'h10030000, 32'h00001003, 32'h00000010, 32'h00001003, 2'b00, 2'b01, 1'bx, 1'b1, 2'b01, 1'b0, 2'b10};
#999 {sound_wr, lights_wr, smem_readdata, dmem_readdata, keyb_char, accel_val, cpu_addr, cpu_readdata, cpu_writedata} <= {1'b0, 1'b0, 32'h00000000, 32'h00000000, 32'h0000001c, 32'h01ea01ea, 32'h10030000, 32'h0000001c, 32'h10010000};

join
end

endmodule